module store_sm (
    start,
    clear,
    clock,
    tready,
    done_,
    tvalid,
    rd_addr,
    rd_en,
    block
);

    input start;
    input clear;
    input clock;
    input tready;
    output done_;
    output tvalid;
    output [5:0] rd_addr;
    output [3:0] rd_en;
    output [1:0] block;

    /* signal declarations */
    wire _45;
    wire _43;
    wire _44;
    wire _41;
    wire _42;
    wire _39;
    wire [1:0] _24;
    wire _38;
    wire _40;
    wire [3:0] _46;
    wire _33;
    wire _31;
    wire _34;
    wire _29;
    wire _35;
    wire _2;
    wire [1:0] _36;
    wire [3:0] _37;
    wire [3:0] _47;
    wire [7:0] _23;
    wire [5:0] _48;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _64;
    wire gnd = 1'b0;
    wire _56;
    wire _57;
    wire _50;
    wire _58;
    wire _49;
    wire _65;
    wire _5;
    reg _53;
    wire [1:0] _26 = 2'b00;
    wire [1:0] _25 = 2'b00;
    wire _8;
    wire [1:0] _94;
    wire [3:0] _62 = 4'b1000;
    wire [3:0] _60 = 4'b0000;
    wire [3:0] _59 = 4'b0000;
    wire [3:0] _72 = 4'b0000;
    wire [3:0] _69 = 4'b0001;
    wire [3:0] _70;
    wire _68;
    wire [3:0] _71;
    wire _67;
    wire [3:0] _73;
    wire [3:0] _9;
    reg [3:0] _61;
    wire _63;
    wire [1:0] _92;
    wire [8:0] _54 = 9'b100001000;
    wire vdd = 1'b1;
    wire [8:0] _20 = 9'b000000000;
    wire _11;
    wire [8:0] _19 = 9'b000000000;
    wire _13;
    wire [8:0] _84 = 9'b000000000;
    wire [8:0] _79 = 9'b000000000;
    wire [8:0] _77 = 9'b000000001;
    wire [8:0] _78;
    wire [8:0] _80;
    wire [8:0] _81;
    wire _76;
    wire [8:0] _82;
    wire _75;
    wire [8:0] _83;
    wire _74;
    wire [8:0] _85;
    wire [8:0] _14;
    reg [8:0] _22;
    wire _55;
    wire [1:0] _89;
    wire _16;
    wire [1:0] _90;
    wire [1:0] _30 = 2'b10;
    wire _88;
    wire [1:0] _91;
    wire [1:0] _28 = 2'b01;
    wire _87;
    wire [1:0] _93;
    wire _86;
    wire [1:0] _95;
    wire [1:0] _17;
    reg [1:0] _27;
    wire [1:0] _66 = 2'b00;
    wire _96;

    /* logic */
    assign _45 = _43 & _41;
    assign _43 = ~ _38;
    assign _44 = _43 & _39;
    assign _41 = ~ _39;
    assign _42 = _38 & _41;
    assign _39 = _24[0:0];
    assign _24 = _23[1:0];
    assign _38 = _24[1:1];
    assign _40 = _38 & _39;
    assign _46 = { _40, _42, _44, _45 };
    assign _33 = _16 ? vdd : gnd;
    assign _31 = _27 == _30;
    assign _34 = _31 ? _33 : gnd;
    assign _29 = _27 == _28;
    assign _35 = _29 ? vdd : _34;
    assign _2 = _35;
    assign _36 = { _2, _2 };
    assign _37 = { _36, _36 };
    assign _47 = _37 & _46;
    assign _23 = _22[7:0];
    assign _48 = _23[7:2];
    assign _64 = _63 ? vdd : _53;
    assign _56 = _55 ? gnd : _53;
    assign _57 = _16 ? _56 : _53;
    assign _50 = _27 == _30;
    assign _58 = _50 ? _57 : _53;
    assign _49 = _27 == _28;
    assign _65 = _49 ? _64 : _58;
    assign _5 = _65;
    always @(posedge _13) begin
        if (_11)
            _53 <= _52;
        else
            _53 <= _5;
    end
    assign _8 = start;
    assign _94 = _8 ? _28 : _27;
    assign _70 = _61 + _69;
    assign _68 = _27 == _28;
    assign _71 = _68 ? _70 : _61;
    assign _67 = _27 == _66;
    assign _73 = _67 ? _72 : _71;
    assign _9 = _73;
    always @(posedge _13) begin
        if (_11)
            _61 <= _60;
        else
            _61 <= _9;
    end
    assign _63 = _61 == _62;
    assign _92 = _63 ? _30 : _27;
    assign _11 = clear;
    assign _13 = clock;
    assign _78 = _22 + _77;
    assign _80 = _55 ? _79 : _78;
    assign _81 = _16 ? _80 : _22;
    assign _76 = _27 == _30;
    assign _82 = _76 ? _81 : _22;
    assign _75 = _27 == _28;
    assign _83 = _75 ? _78 : _82;
    assign _74 = _27 == _66;
    assign _85 = _74 ? _84 : _83;
    assign _14 = _85;
    always @(posedge _13) begin
        if (_11)
            _22 <= _20;
        else
            _22 <= _14;
    end
    assign _55 = _22 == _54;
    assign _89 = _55 ? _66 : _27;
    assign _16 = tready;
    assign _90 = _16 ? _89 : _27;
    assign _88 = _27 == _30;
    assign _91 = _88 ? _90 : _27;
    assign _87 = _27 == _28;
    assign _93 = _87 ? _92 : _91;
    assign _86 = _27 == _66;
    assign _95 = _86 ? _94 : _93;
    assign _17 = _95;
    always @(posedge _13) begin
        if (_11)
            _27 <= _26;
        else
            _27 <= _17;
    end
    assign _96 = _66 == _27;

    /* aliases */

    /* output assignments */
    assign done_ = _96;
    assign tvalid = _53;
    assign rd_addr = _48;
    assign rd_en = _47;
    assign block = _24;

endmodule
module controller (
    start,
    clear,
    clock,
    cores_done,
    output_done,
    input_done,
    done_,
    start_input,
    start_output,
    start_cores,
    first_iter,
    flip
);

    input start;
    input clear;
    input clock;
    input cores_done;
    input output_done;
    input input_done;
    output done_;
    output start_input;
    output start_output;
    output start_cores;
    output first_iter;
    output flip;

    /* signal declarations */
    wire _25;
    wire _35 = 1'b1;
    wire _36;
    wire _31;
    wire _37;
    wire _2;
    wire _51;
    wire _48;
    wire _49;
    wire _40;
    wire _50;
    wire _38;
    wire _52;
    wire START_CORES;
    wire _58;
    wire _59;
    wire _56;
    wire _55;
    wire _57;
    wire _53;
    wire _60;
    wire START_OUTPUT;
    wire _70;
    wire _68;
    wire _65;
    wire _66;
    wire gnd = 1'b0;
    wire _64;
    wire _67;
    wire _63;
    wire _69;
    wire _62;
    wire _71;
    wire START_INPUT;
    wire [2:0] _27 = 3'b000;
    wire [2:0] _26 = 3'b000;
    wire _11;
    wire [2:0] _94;
    wire [2:0] _92;
    wire _46 = 1'b0;
    wire _44 = 1'b1;
    wire vdd = 1'b1;
    wire _42 = 1'b0;
    wire _13;
    wire _41 = 1'b0;
    wire _15;
    wire _76 = 1'b1;
    wire _77;
    wire _74;
    wire _73;
    wire _75;
    wire _72;
    wire _78;
    wire _16;
    reg ITERATION;
    wire _45;
    wire _47;
    wire [2:0] _89;
    wire [2:0] _90;
    wire [2:0] _87;
    wire _18;
    wire _20;
    wire _22;
    wire _33;
    wire _34;
    wire [2:0] _85;
    wire [2:0] _83 = 3'b100;
    wire _84;
    wire [2:0] _86;
    wire [2:0] _54 = 3'b011;
    wire _82;
    wire [2:0] _88;
    wire [2:0] _39 = 3'b010;
    wire _81;
    wire [2:0] _91;
    wire [2:0] _30 = 3'b001;
    wire _80;
    wire [2:0] _93;
    wire _79;
    wire [2:0] _95;
    wire [2:0] _23;
    reg [2:0] STATE;
    wire [2:0] _61 = 3'b000;
    wire _96;

    /* logic */
    assign _25 = START_CORES | START_OUTPUT;
    assign _36 = _34 ? _35 : gnd;
    assign _31 = STATE == _30;
    assign _37 = _31 ? _36 : gnd;
    assign _2 = _37;
    assign _51 = _34 ? vdd : gnd;
    assign _48 = _47 ? vdd : vdd;
    assign _49 = _34 ? _48 : gnd;
    assign _40 = STATE == _39;
    assign _50 = _40 ? _49 : gnd;
    assign _38 = STATE == _30;
    assign _52 = _38 ? _51 : _50;
    assign START_CORES = _52;
    assign _58 = _47 ? vdd : vdd;
    assign _59 = _34 ? _58 : gnd;
    assign _56 = _34 ? vdd : gnd;
    assign _55 = STATE == _54;
    assign _57 = _55 ? _56 : gnd;
    assign _53 = STATE == _39;
    assign _60 = _53 ? _59 : _57;
    assign START_OUTPUT = _60;
    assign _70 = _11 ? vdd : gnd;
    assign _68 = _34 ? vdd : gnd;
    assign _65 = _47 ? gnd : vdd;
    assign _66 = _34 ? _65 : gnd;
    assign _64 = STATE == _39;
    assign _67 = _64 ? _66 : gnd;
    assign _63 = STATE == _30;
    assign _69 = _63 ? _68 : _67;
    assign _62 = STATE == _61;
    assign _71 = _62 ? _70 : _69;
    assign START_INPUT = _71;
    assign _11 = start;
    assign _94 = _11 ? _30 : STATE;
    assign _92 = _34 ? _39 : STATE;
    assign _13 = clear;
    assign _15 = clock;
    assign _77 = _34 ? _76 : ITERATION;
    assign _74 = _34 ? _45 : ITERATION;
    assign _73 = STATE == _39;
    assign _75 = _73 ? _74 : ITERATION;
    assign _72 = STATE == _30;
    assign _78 = _72 ? _77 : _75;
    assign _16 = _78;
    always @(posedge _15) begin
        if (_13)
            ITERATION <= _42;
        else
            ITERATION <= _16;
    end
    assign _45 = ITERATION + _44;
    assign _47 = _45 == _46;
    assign _89 = _47 ? _54 : STATE;
    assign _90 = _34 ? _89 : STATE;
    assign _87 = _34 ? _83 : STATE;
    assign _18 = cores_done;
    assign _20 = output_done;
    assign _22 = input_done;
    assign _33 = _22 & _20;
    assign _34 = _33 & _18;
    assign _85 = _34 ? _61 : STATE;
    assign _84 = STATE == _83;
    assign _86 = _84 ? _85 : STATE;
    assign _82 = STATE == _54;
    assign _88 = _82 ? _87 : _86;
    assign _81 = STATE == _39;
    assign _91 = _81 ? _90 : _88;
    assign _80 = STATE == _30;
    assign _93 = _80 ? _92 : _91;
    assign _79 = STATE == _61;
    assign _95 = _79 ? _94 : _93;
    assign _23 = _95;
    always @(posedge _15) begin
        if (_13)
            STATE <= _27;
        else
            STATE <= _23;
    end
    assign _96 = _61 == STATE;

    /* aliases */

    /* output assignments */
    assign done_ = _96;
    assign start_input = START_INPUT;
    assign start_output = START_OUTPUT;
    assign start_cores = START_CORES;
    assign first_iter = _2;
    assign flip = _25;

endmodule
module load_sm (
    first_4step_pass,
    start,
    tvalid,
    clear,
    clock,
    done_,
    tready,
    wr_addr,
    wr_en
);

    input first_4step_pass;
    input start;
    input tvalid;
    input clear;
    input clock;
    output done_;
    output tready;
    output [5:0] wr_addr;
    output [3:0] wr_en;

    /* signal declarations */
    wire _40;
    wire _38;
    wire _39;
    wire _36;
    wire _37;
    wire _34;
    wire [1:0] _31;
    wire [1:0] _30;
    wire [1:0] _32;
    wire _33;
    wire _35;
    wire [3:0] _41;
    wire _24;
    wire [1:0] _25;
    wire [3:0] _26;
    wire [3:0] _42;
    wire [5:0] _44;
    wire [5:0] _43;
    wire _3;
    wire [5:0] _45;
    wire _23;
    wire [1:0] _20 = 2'b00;
    wire [1:0] _19 = 2'b00;
    wire _7;
    wire [1:0] _78;
    wire [7:0] _73 = 8'b00000000;
    wire [7:0] _49 = 8'b00000001;
    wire [7:0] _28 = 8'b00000000;
    wire [7:0] _27 = 8'b00000000;
    wire [7:0] _53 = 8'b00000000;
    wire [7:0] _51;
    wire _48;
    wire [7:0] _52;
    wire _47;
    wire [7:0] _54;
    wire [7:0] _8;
    reg [7:0] _29;
    wire [7:0] _50;
    wire _74;
    wire [1:0] _75;
    wire _10;
    wire [1:0] _76;
    wire _69 = 1'b1;
    wire vdd = 1'b1;
    wire _59 = 1'b0;
    wire _12;
    wire _58 = 1'b0;
    wire _14;
    wire _64 = 1'b0;
    wire _61 = 1'b1;
    wire _62;
    wire _57;
    wire _63;
    wire _55;
    wire _65;
    wire _15;
    reg _60;
    wire _70;
    wire [1:0] _71;
    wire [1:0] _56 = 2'b10;
    wire _68;
    wire [1:0] _72;
    wire [1:0] _18 = 2'b01;
    wire _67;
    wire [1:0] _77;
    wire _66;
    wire [1:0] _79;
    wire [1:0] _16;
    reg [1:0] _22;
    wire [1:0] _46 = 2'b00;
    wire _80;

    /* logic */
    assign _40 = _38 & _36;
    assign _38 = ~ _33;
    assign _39 = _38 & _34;
    assign _36 = ~ _34;
    assign _37 = _33 & _36;
    assign _34 = _32[0:0];
    assign _31 = _29[1:0];
    assign _30 = _29[7:6];
    assign _32 = _3 ? _31 : _30;
    assign _33 = _32[1:1];
    assign _35 = _33 & _34;
    assign _41 = { _35, _37, _39, _40 };
    assign _24 = _23 & _10;
    assign _25 = { _24, _24 };
    assign _26 = { _25, _25 };
    assign _42 = _26 & _41;
    assign _44 = _29[7:2];
    assign _43 = _29[5:0];
    assign _3 = first_4step_pass;
    assign _45 = _3 ? _44 : _43;
    assign _23 = _18 == _22;
    assign _7 = start;
    assign _78 = _7 ? _18 : _22;
    assign _51 = _10 ? _50 : _29;
    assign _48 = _22 == _18;
    assign _52 = _48 ? _51 : _29;
    assign _47 = _22 == _46;
    assign _54 = _47 ? _53 : _52;
    assign _8 = _54;
    always @(posedge _14) begin
        if (_12)
            _29 <= _28;
        else
            _29 <= _8;
    end
    assign _50 = _29 + _49;
    assign _74 = _50 == _73;
    assign _75 = _74 ? _56 : _22;
    assign _10 = tvalid;
    assign _76 = _10 ? _75 : _22;
    assign _12 = clear;
    assign _14 = clock;
    assign _62 = _60 + _61;
    assign _57 = _22 == _56;
    assign _63 = _57 ? _62 : _60;
    assign _55 = _22 == _46;
    assign _65 = _55 ? _64 : _63;
    assign _15 = _65;
    always @(posedge _14) begin
        if (_12)
            _60 <= _59;
        else
            _60 <= _15;
    end
    assign _70 = _60 == _69;
    assign _71 = _70 ? _46 : _22;
    assign _68 = _22 == _56;
    assign _72 = _68 ? _71 : _22;
    assign _67 = _22 == _18;
    assign _77 = _67 ? _76 : _72;
    assign _66 = _22 == _46;
    assign _79 = _66 ? _78 : _77;
    assign _16 = _79;
    always @(posedge _14) begin
        if (_12)
            _22 <= _20;
        else
            _22 <= _16;
    end
    assign _80 = _46 == _22;

    /* aliases */

    /* output assignments */
    assign done_ = _80;
    assign tready = _23;
    assign wr_addr = _45;
    assign wr_en = _42;

endmodule
module ctrl (
    first_4step_pass,
    start,
    clear,
    clock,
    first_iter,
    done_,
    i,
    j,
    k,
    m,
    addr1,
    addr2,
    omegas0,
    omegas1,
    omegas2,
    omegas3,
    omegas4,
    omegas5,
    omegas6,
    start_twiddles,
    first_stage,
    last_stage,
    twiddle_stage,
    valid,
    index,
    read_write_enable,
    flip
);

    input first_4step_pass;
    input start;
    input clear;
    input clock;
    input first_iter;
    output done_;
    output [2:0] i;
    output [5:0] j;
    output [5:0] k;
    output [5:0] m;
    output [5:0] addr1;
    output [5:0] addr2;
    output [63:0] omegas0;
    output [63:0] omegas1;
    output [63:0] omegas2;
    output [63:0] omegas3;
    output [63:0] omegas4;
    output [63:0] omegas5;
    output [63:0] omegas6;
    output start_twiddles;
    output first_stage;
    output last_stage;
    output twiddle_stage;
    output valid;
    output [3:0] index;
    output read_write_enable;
    output flip;

    /* signal declarations */
    wire _59;
    wire _52;
    wire _60;
    wire _1;
    wire _64;
    wire _65;
    wire _62;
    wire _66;
    wire _3;
    wire _73 = 1'b0;
    wire _72 = 1'b0;
    wire _92 = 1'b0;
    wire _93;
    wire _89 = 1'b1;
    wire _90;
    wire _81 = 1'b0;
    wire _79 = 1'b0;
    wire [3:0] _77 = 4'b0110;
    wire _78;
    wire _80;
    wire _82;
    wire _71;
    wire _83;
    wire _69;
    wire _91;
    wire _68;
    wire _94;
    wire _6;
    reg _74;
    wire _100 = 1'b0;
    wire _99 = 1'b0;
    wire _120 = 1'b0;
    wire _121;
    wire _115 = 1'b1;
    wire _116;
    wire _117;
    wire _118;
    wire _105 = 1'b0;
    wire _106;
    wire _102 = 1'b0;
    wire _103;
    wire _98;
    wire _104;
    wire _97;
    wire _107;
    wire _96;
    wire _119;
    wire _95;
    wire _122;
    wire _8;
    reg _101;
    wire _127 = 1'b0;
    wire _126 = 1'b0;
    wire _141 = 1'b0;
    wire _142;
    wire _136 = 1'b1;
    wire _135 = 1'b0;
    wire _137;
    wire _133;
    wire [2:0] _131 = 3'b101;
    wire _132;
    wire _134;
    wire _138;
    wire _139;
    wire gnd = 1'b0;
    wire _129;
    wire _125;
    wire _130;
    wire _124;
    wire _140;
    wire _123;
    wire _143;
    wire _10;
    reg _128;
    wire _147 = 1'b0;
    wire _146 = 1'b0;
    wire _152 = 1'b1;
    wire _153;
    wire _149 = 1'b0;
    wire _150;
    wire _145;
    wire _151;
    wire _144;
    wire _154;
    wire _12;
    reg _148;
    wire _188 = 1'b0;
    wire _187 = 1'b0;
    wire _184 = 1'b1;
    wire _185;
    wire _180 = 1'b1;
    wire _181;
    wire _182;
    wire _159 = 1'b1;
    wire _160;
    wire _158 = 1'b0;
    wire _157;
    wire _161;
    wire _156;
    wire _183;
    wire _155;
    wire _186;
    wire _14;
    reg _189;
    wire [63:0] _195 = 64'b0000000000000001111111111111111111111111111111100000000000000000;
    wire [63:0] _194 = 64'b1111111111111111111111111111101100000000000000000000000000000101;
    wire [63:0] _193 = 64'b1111111111111111111111111110111100000000000000000000000000000001;
    wire [63:0] _192 = 64'b0000000000000000000000001111111111111111111111111111111100000000;
    wire [63:0] _191 = 64'b1111111111111110111111111111111100000000000000000000000000000001;
    wire [63:0] _190 = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    reg [63:0] _196;
    wire [63:0] _202 = 64'b0000000000000000000001000000000000000000000000000000000000000000;
    wire [63:0] _201 = 64'b0000000000001111111111111111111111111111111100000000000000000000;
    wire [63:0] _200 = 64'b1111111111111111111111101111111100000000000000000000000100000001;
    wire [63:0] _199 = 64'b1111111111111110111111111111111100000000000000000000000000000001;
    wire [63:0] _198 = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [63:0] _197 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    reg [63:0] _203;
    wire [63:0] _209 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    wire [63:0] _208 = 64'b0000000000000000000000000000000000000000000000000000000001000000;
    wire [63:0] _207 = 64'b0000000000000000000000000000000000000000000000000001000000000000;
    wire [63:0] _206 = 64'b0000000000000000000000000000000000000001000000000000000000000000;
    wire [63:0] _205 = 64'b0000000000000001000000000000000000000000000000000000000000000000;
    wire [63:0] _204 = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    reg [63:0] _210;
    wire [63:0] _216 = 64'b1110111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _215 = 64'b1111111111111111111111111111111011111111000000000000000000000001;
    wire [63:0] _214 = 64'b0000000000000001000000000000000000000000000000000000000000000000;
    wire [63:0] _213 = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _211 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    reg [63:0] _217;
    wire [63:0] _223 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _222 = 64'b0000000000000000000001000000000000000000000000000000000000000000;
    wire [63:0] _221 = 64'b0000000000001111111111111111111111111111111100000000000000000000;
    wire [63:0] _220 = 64'b1111111111111111111111101111111100000000000000000000000100000001;
    wire [63:0] _219 = 64'b1111111111111110111111111111111100000000000000000000000000000001;
    wire [63:0] _218 = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    reg [63:0] _224;
    wire [63:0] _230 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _229 = 64'b1110111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _228 = 64'b1111111111111111111111111111111011111111000000000000000000000001;
    wire [63:0] _227 = 64'b0000000000000001000000000000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [63:0] _225 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    reg [63:0] _231;
    wire [63:0] _237 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _235 = 64'b1110111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _234 = 64'b1111111111111111111111111111111011111111000000000000000000000001;
    wire [63:0] _233 = 64'b0000000000000001000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    reg [63:0] _238;
    wire [5:0] _243 = 6'b000000;
    wire [5:0] _242 = 6'b000000;
    wire [5:0] _252 = 6'b000000;
    wire [5:0] _253;
    wire [5:0] _249;
    wire [5:0] _247 = 6'b000001;
    wire [5:0] _248;
    wire [5:0] _250;
    wire [5:0] _245;
    wire _241;
    wire [5:0] _246;
    wire _240;
    wire [5:0] _251;
    wire _239;
    wire [5:0] _254;
    wire [5:0] _24;
    reg [5:0] _244;
    wire _344 = 1'b0;
    wire _354 = 1'b0;
    wire _355;
    wire _349 = 1'b1;
    wire _350;
    wire _351;
    wire _352;
    wire _346 = 1'b1;
    wire _347;
    wire _343;
    wire _348;
    wire _342;
    wire _353;
    wire [2:0] _48 = 3'b000;
    wire [2:0] _47 = 3'b000;
    wire [2:0] _339;
    wire [2:0] _336;
    wire [2:0] _337;
    wire [2:0] _332;
    wire [2:0] _333;
    wire [2:0] _334;
    wire [5:0] _87 = 6'b111111;
    wire [5:0] _85 = 6'b000000;
    wire [5:0] _84 = 6'b000000;
    wire [5:0] _312 = 6'b000001;
    wire [5:0] _313;
    wire [5:0] _308;
    wire [5:0] _309;
    wire [5:0] _310;
    wire [5:0] _303 = 6'b000000;
    wire _31;
    wire [5:0] _304;
    wire [5:0] _172 = 6'b000000;
    wire [5:0] _171 = 6'b000000;
    wire [5:0] _283 = 6'b000000;
    wire [5:0] _284;
    wire [5:0] _280;
    wire [5:0] _168 = 6'b000000;
    wire [5:0] _167 = 6'b000000;
    wire [5:0] _259 = 6'b000001;
    wire [5:0] _260;
    wire _175 = 1'b0;
    wire [4:0] _174;
    wire [5:0] _176;
    wire [5:0] _257;
    wire _256;
    wire [5:0] _258;
    wire _255;
    wire [5:0] _261;
    wire [5:0] _32;
    reg [5:0] m_0;
    wire [5:0] _165 = 6'b000001;
    wire [5:0] _163 = 6'b000000;
    wire [5:0] _162 = 6'b000000;
    wire [5:0] _272 = 6'b000000;
    wire [5:0] _273;
    wire [5:0] _268 = 6'b000000;
    wire [5:0] _178 = 6'b000000;
    wire _179;
    wire [5:0] _269;
    wire [5:0] _270;
    wire [5:0] _265 = 6'b000000;
    wire [5:0] _266;
    wire _264;
    wire [5:0] _267;
    wire _263;
    wire [5:0] _271;
    wire _262;
    wire [5:0] _274;
    wire [5:0] _33;
    reg [5:0] j_0;
    wire [5:0] _166;
    wire _170;
    wire [5:0] _281;
    wire [5:0] _278;
    wire _277;
    wire [5:0] _279;
    wire _276;
    wire [5:0] _282;
    wire _275;
    wire [5:0] _285;
    wire [5:0] _34;
    reg [5:0] k_0;
    wire [5:0] _177;
    wire [5:0] _302;
    wire [2:0] _113 = 3'b110;
    wire [2:0] _111 = 3'b001;
    wire [2:0] _109 = 3'b000;
    wire [2:0] _108 = 3'b000;
    wire [2:0] _290 = 3'b000;
    wire _36;
    wire [2:0] _291;
    wire [2:0] _288;
    wire _287;
    wire [2:0] _289;
    wire _286;
    wire [2:0] _292;
    wire [2:0] _37;
    reg [2:0] i_0;
    wire [2:0] _112;
    wire _114;
    wire [5:0] _305;
    wire [5:0] _306;
    wire [5:0] _299 = 6'b000000;
    wire [5:0] _297 = 6'b000001;
    wire [5:0] _298;
    wire [5:0] _300;
    wire _296;
    wire [5:0] _301;
    wire _295;
    wire [5:0] _307;
    wire _294;
    wire [5:0] _311;
    wire _293;
    wire [5:0] _314;
    wire [5:0] _38;
    reg [5:0] _86;
    wire _88;
    wire [2:0] _330;
    wire [3:0] _75 = 4'b1000;
    wire vdd = 1'b1;
    wire [3:0] _55 = 4'b0000;
    wire _40;
    wire [3:0] _54 = 4'b0000;
    wire _42;
    wire [3:0] _320 = 4'b0000;
    wire [3:0] _57 = 4'b1000;
    wire _58;
    wire [3:0] _321;
    wire [3:0] _317 = 4'b0001;
    wire [3:0] _318;
    wire _316;
    wire [3:0] _319;
    wire _315;
    wire [3:0] _322;
    wire [3:0] _43;
    reg [3:0] _56;
    wire _76;
    wire [2:0] _328;
    wire [2:0] _70 = 3'b100;
    wire _327;
    wire [2:0] _329;
    wire [2:0] _63 = 3'b011;
    wire _326;
    wire [2:0] _331;
    wire [2:0] _51 = 3'b010;
    wire _325;
    wire [2:0] _335;
    wire [2:0] _61 = 3'b001;
    wire _324;
    wire [2:0] _338;
    wire [2:0] _67 = 3'b000;
    wire _323;
    wire [2:0] _340;
    wire [2:0] _44;
    reg [2:0] STATE;
    wire _341;
    wire _356;
    wire _45;
    reg _345;

    /* logic */
    assign _59 = _58 ? vdd : gnd;
    assign _52 = STATE == _51;
    assign _60 = _52 ? _59 : gnd;
    assign _1 = _60;
    assign _64 = STATE == _63;
    assign _65 = _64 ? vdd : gnd;
    assign _62 = STATE == _61;
    assign _66 = _62 ? vdd : _65;
    assign _3 = _66;
    assign _93 = _36 ? _92 : _74;
    assign _90 = _88 ? _89 : _74;
    assign _78 = _56 == _77;
    assign _80 = _78 ? _79 : _74;
    assign _82 = _76 ? _81 : _80;
    assign _71 = STATE == _70;
    assign _83 = _71 ? _82 : _74;
    assign _69 = STATE == _63;
    assign _91 = _69 ? _90 : _83;
    assign _68 = STATE == _67;
    assign _94 = _68 ? _93 : _91;
    assign _6 = _94;
    always @(posedge _42) begin
        if (_40)
            _74 <= _73;
        else
            _74 <= _6;
    end
    assign _121 = _36 ? _120 : _101;
    assign _116 = _31 ? _115 : _101;
    assign _117 = _114 ? _116 : _101;
    assign _118 = _58 ? _117 : _101;
    assign _106 = _88 ? _105 : _101;
    assign _103 = _76 ? _102 : _101;
    assign _98 = STATE == _70;
    assign _104 = _98 ? _103 : _101;
    assign _97 = STATE == _63;
    assign _107 = _97 ? _106 : _104;
    assign _96 = STATE == _51;
    assign _119 = _96 ? _118 : _107;
    assign _95 = STATE == _67;
    assign _122 = _95 ? _121 : _119;
    assign _8 = _122;
    always @(posedge _42) begin
        if (_40)
            _101 <= _100;
        else
            _101 <= _8;
    end
    assign _142 = _36 ? _141 : _128;
    assign _137 = _31 ? _136 : _135;
    assign _133 = ~ _31;
    assign _132 = _112 == _131;
    assign _134 = _132 ? _133 : _128;
    assign _138 = _114 ? _137 : _134;
    assign _139 = _58 ? _138 : _128;
    assign _129 = _76 ? gnd : _128;
    assign _125 = STATE == _70;
    assign _130 = _125 ? _129 : _128;
    assign _124 = STATE == _51;
    assign _140 = _124 ? _139 : _130;
    assign _123 = STATE == _67;
    assign _143 = _123 ? _142 : _140;
    assign _10 = _143;
    always @(posedge _42) begin
        if (_40)
            _128 <= _127;
        else
            _128 <= _10;
    end
    assign _153 = _36 ? _152 : _148;
    assign _150 = _58 ? _149 : _148;
    assign _145 = STATE == _51;
    assign _151 = _145 ? _150 : _148;
    assign _144 = STATE == _67;
    assign _154 = _144 ? _153 : _151;
    assign _12 = _154;
    always @(posedge _42) begin
        if (_40)
            _148 <= _147;
        else
            _148 <= _12;
    end
    assign _185 = _36 ? _184 : _158;
    assign _181 = _179 ? _158 : _180;
    assign _182 = _170 ? _181 : _158;
    assign _160 = _58 ? _159 : _158;
    assign _157 = STATE == _51;
    assign _161 = _157 ? _160 : _158;
    assign _156 = STATE == _61;
    assign _183 = _156 ? _182 : _161;
    assign _155 = STATE == _67;
    assign _186 = _155 ? _185 : _183;
    assign _14 = _186;
    always @(posedge _42) begin
        if (_40)
            _189 <= _188;
        else
            _189 <= _14;
    end
    always @* begin
        case (i_0)
        0: _196 <= _190;
        1: _196 <= _191;
        2: _196 <= _192;
        3: _196 <= _193;
        4: _196 <= _194;
        default: _196 <= _195;
        endcase
    end
    always @* begin
        case (i_0)
        0: _203 <= _197;
        1: _203 <= _198;
        2: _203 <= _199;
        3: _203 <= _200;
        4: _203 <= _201;
        default: _203 <= _202;
        endcase
    end
    always @* begin
        case (i_0)
        0: _210 <= _204;
        1: _210 <= _205;
        2: _210 <= _206;
        3: _210 <= _207;
        4: _210 <= _208;
        default: _210 <= _209;
        endcase
    end
    always @* begin
        case (i_0)
        0: _217 <= _211;
        1: _217 <= _212;
        2: _217 <= _213;
        3: _217 <= _214;
        4: _217 <= _215;
        default: _217 <= _216;
        endcase
    end
    always @* begin
        case (i_0)
        0: _224 <= _218;
        1: _224 <= _219;
        2: _224 <= _220;
        3: _224 <= _221;
        4: _224 <= _222;
        default: _224 <= _223;
        endcase
    end
    always @* begin
        case (i_0)
        0: _231 <= _225;
        1: _231 <= _226;
        2: _231 <= _227;
        3: _231 <= _228;
        4: _231 <= _229;
        default: _231 <= _230;
        endcase
    end
    always @* begin
        case (i_0)
        0: _238 <= _232;
        1: _238 <= _233;
        2: _238 <= _234;
        3: _238 <= _235;
        4: _238 <= _236;
        default: _238 <= _237;
        endcase
    end
    assign _253 = _36 ? _252 : _244;
    assign _249 = _179 ? _248 : _177;
    assign _248 = _244 + _247;
    assign _250 = _170 ? _249 : _248;
    assign _245 = _58 ? _177 : _244;
    assign _241 = STATE == _51;
    assign _246 = _241 ? _245 : _244;
    assign _240 = STATE == _61;
    assign _251 = _240 ? _250 : _246;
    assign _239 = STATE == _67;
    assign _254 = _239 ? _253 : _251;
    assign _24 = _254;
    always @(posedge _42) begin
        if (_40)
            _244 <= _243;
        else
            _244 <= _24;
    end
    assign _355 = _36 ? _354 : _345;
    assign _350 = _31 ? _345 : _349;
    assign _351 = _114 ? _350 : _345;
    assign _352 = _58 ? _351 : _345;
    assign _347 = _76 ? _346 : _345;
    assign _343 = STATE == _70;
    assign _348 = _343 ? _347 : _345;
    assign _342 = STATE == _51;
    assign _353 = _342 ? _352 : _348;
    assign _339 = _36 ? _61 : STATE;
    assign _336 = _179 ? _51 : STATE;
    assign _337 = _170 ? _336 : STATE;
    assign _332 = _31 ? _63 : _67;
    assign _333 = _114 ? _332 : _61;
    assign _334 = _58 ? _333 : STATE;
    assign _313 = _36 ? _312 : _86;
    assign _308 = _177 + m_0;
    assign _309 = _179 ? _298 : _308;
    assign _310 = _170 ? _309 : _298;
    assign _31 = first_4step_pass;
    assign _304 = _31 ? _303 : _302;
    assign _284 = _36 ? _283 : k_0;
    assign _280 = _179 ? k_0 : _177;
    assign _260 = _36 ? _259 : m_0;
    assign _174 = m_0[4:0];
    assign _176 = { _174, _175 };
    assign _257 = _58 ? _176 : m_0;
    assign _256 = STATE == _51;
    assign _258 = _256 ? _257 : m_0;
    assign _255 = STATE == _67;
    assign _261 = _255 ? _260 : _258;
    assign _32 = _261;
    always @(posedge _42) begin
        if (_40)
            m_0 <= _168;
        else
            m_0 <= _32;
    end
    assign _273 = _36 ? _272 : j_0;
    assign _179 = _177 == _178;
    assign _269 = _179 ? _166 : _268;
    assign _270 = _170 ? _269 : _166;
    assign _266 = _58 ? _265 : j_0;
    assign _264 = STATE == _51;
    assign _267 = _264 ? _266 : j_0;
    assign _263 = STATE == _61;
    assign _271 = _263 ? _270 : _267;
    assign _262 = STATE == _67;
    assign _274 = _262 ? _273 : _271;
    assign _33 = _274;
    always @(posedge _42) begin
        if (_40)
            j_0 <= _163;
        else
            j_0 <= _33;
    end
    assign _166 = j_0 + _165;
    assign _170 = _166 == m_0;
    assign _281 = _170 ? _280 : k_0;
    assign _278 = _58 ? _177 : k_0;
    assign _277 = STATE == _51;
    assign _279 = _277 ? _278 : k_0;
    assign _276 = STATE == _61;
    assign _282 = _276 ? _281 : _279;
    assign _275 = STATE == _67;
    assign _285 = _275 ? _284 : _282;
    assign _34 = _285;
    always @(posedge _42) begin
        if (_40)
            k_0 <= _172;
        else
            k_0 <= _34;
    end
    assign _177 = k_0 + _176;
    assign _302 = _177 + _176;
    assign _36 = start;
    assign _291 = _36 ? _290 : i_0;
    assign _288 = _58 ? _112 : i_0;
    assign _287 = STATE == _51;
    assign _289 = _287 ? _288 : i_0;
    assign _286 = STATE == _67;
    assign _292 = _286 ? _291 : _289;
    assign _37 = _292;
    always @(posedge _42) begin
        if (_40)
            i_0 <= _109;
        else
            i_0 <= _37;
    end
    assign _112 = i_0 + _111;
    assign _114 = _112 == _113;
    assign _305 = _114 ? _304 : _302;
    assign _306 = _58 ? _305 : _86;
    assign _298 = _86 + _297;
    assign _300 = _88 ? _299 : _298;
    assign _296 = STATE == _63;
    assign _301 = _296 ? _300 : _86;
    assign _295 = STATE == _51;
    assign _307 = _295 ? _306 : _301;
    assign _294 = STATE == _61;
    assign _311 = _294 ? _310 : _307;
    assign _293 = STATE == _67;
    assign _314 = _293 ? _313 : _311;
    assign _38 = _314;
    always @(posedge _42) begin
        if (_40)
            _86 <= _85;
        else
            _86 <= _38;
    end
    assign _88 = _86 == _87;
    assign _330 = _88 ? _70 : STATE;
    assign _40 = clear;
    assign _42 = clock;
    assign _58 = _56 == _57;
    assign _321 = _58 ? _320 : _318;
    assign _318 = _56 + _317;
    assign _316 = STATE == _70;
    assign _319 = _316 ? _318 : _56;
    assign _315 = STATE == _51;
    assign _322 = _315 ? _321 : _319;
    assign _43 = _322;
    always @(posedge _42) begin
        if (_40)
            _56 <= _55;
        else
            _56 <= _43;
    end
    assign _76 = _56 == _75;
    assign _328 = _76 ? _67 : STATE;
    assign _327 = STATE == _70;
    assign _329 = _327 ? _328 : STATE;
    assign _326 = STATE == _63;
    assign _331 = _326 ? _330 : _329;
    assign _325 = STATE == _51;
    assign _335 = _325 ? _334 : _331;
    assign _324 = STATE == _61;
    assign _338 = _324 ? _337 : _335;
    assign _323 = STATE == _67;
    assign _340 = _323 ? _339 : _338;
    assign _44 = _340;
    always @(posedge _42) begin
        if (_40)
            STATE <= _48;
        else
            STATE <= _44;
    end
    assign _341 = STATE == _67;
    assign _356 = _341 ? _355 : _353;
    assign _45 = _356;
    always @(posedge _42) begin
        if (_40)
            _345 <= vdd;
        else
            _345 <= _45;
    end

    /* aliases */

    /* output assignments */
    assign done_ = _345;
    assign i = i_0;
    assign j = j_0;
    assign k = k_0;
    assign m = m_0;
    assign addr1 = _244;
    assign addr2 = _86;
    assign omegas0 = _238;
    assign omegas1 = _231;
    assign omegas2 = _224;
    assign omegas3 = _217;
    assign omegas4 = _210;
    assign omegas5 = _203;
    assign omegas6 = _196;
    assign start_twiddles = _189;
    assign first_stage = _148;
    assign last_stage = _128;
    assign twiddle_stage = _101;
    assign valid = _74;
    assign index = _56;
    assign read_write_enable = _3;
    assign flip = _1;

endmodule
module twdl (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    clock,
    start_twiddles,
    w
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input clock;
    input start_twiddles;
    output [63:0] w;

    /* signal declarations */
    wire [63:0] _36 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _35 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _87 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _83 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _84;
    wire [64:0] _80 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _77 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _76 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _73 = 33'b000000000000000000000000000000000;
    wire [64:0] _74;
    wire [31:0] _70 = 32'b00000000000000000000000000000000;
    wire [31:0] _69;
    wire [63:0] _71;
    wire [64:0] _72;
    wire [64:0] _75;
    reg [64:0] _78;
    wire [64:0] _67 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _66 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _63 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _61;
    wire [64:0] _62;
    wire [64:0] _64;
    wire [31:0] _57;
    wire [32:0] _56 = 33'b000000000000000000000000000000000;
    wire [64:0] _58;
    wire [127:0] _52 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _51 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _49 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _48 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _46 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _45 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _42 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _41 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _2;
    reg [63:0] _43;
    wire [63:0] _39 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    reg [63:0] _40;
    wire [127:0] _44;
    reg [127:0] _47;
    reg [127:0] _50;
    reg [127:0] _53;
    wire [63:0] _54;
    wire gnd = 1'b0;
    wire [64:0] _55;
    wire [64:0] _59;
    wire _60;
    wire [64:0] _65;
    reg [64:0] _68;
    wire [64:0] _79;
    wire _81;
    wire _82;
    wire [64:0] _85;
    wire [63:0] _86;
    reg [63:0] _89;
    wire [63:0] _4;
    wire [63:0] _6;
    wire [63:0] _8;
    wire [63:0] _10;
    wire [63:0] _12;
    wire [63:0] _14;
    wire vdd = 1'b1;
    wire [2:0] _23 = 3'b000;
    wire [2:0] _22 = 3'b000;
    wire _16;
    wire [2:0] _32 = 3'b000;
    wire [2:0] _29 = 3'b001;
    wire [2:0] _30;
    wire [2:0] _26 = 3'b110;
    wire _27;
    wire _28;
    wire [2:0] _31;
    wire [2:0] _33;
    wire [2:0] _17;
    reg [2:0] _25;
    reg [63:0] _90;
    wire _19;
    wire [63:0] _92;
    wire [63:0] _20;
    reg [63:0] _37;

    /* logic */
    assign _84 = _79 - _83;
    assign _74 = { _73, _69 };
    assign _69 = _53[95:64];
    assign _71 = { _69, _70 };
    assign _72 = { gnd, _71 };
    assign _75 = _72 - _74;
    always @(posedge _16) begin
        _78 <= _75;
    end
    assign _61 = _59[63:0];
    assign _62 = { gnd, _61 };
    assign _64 = _62 - _63;
    assign _57 = _53[127:96];
    assign _58 = { _56, _57 };
    assign _2 = omegas6;
    always @(posedge _16) begin
        _43 <= _2;
    end
    always @(posedge _16) begin
        _40 <= _37;
    end
    assign _44 = _40 * _43;
    always @(posedge _16) begin
        _47 <= _44;
    end
    always @(posedge _16) begin
        _50 <= _47;
    end
    always @(posedge _16) begin
        _53 <= _50;
    end
    assign _54 = _53[63:0];
    assign _55 = { gnd, _54 };
    assign _59 = _55 - _58;
    assign _60 = _59[64:64];
    assign _65 = _60 ? _64 : _59;
    always @(posedge _16) begin
        _68 <= _65;
    end
    assign _79 = _68 + _78;
    assign _81 = _79 < _80;
    assign _82 = ~ _81;
    assign _85 = _82 ? _84 : _79;
    assign _86 = _85[63:0];
    always @(posedge _16) begin
        _89 <= _86;
    end
    assign _4 = omegas5;
    assign _6 = omegas4;
    assign _8 = omegas3;
    assign _10 = omegas2;
    assign _12 = omegas1;
    assign _14 = omegas0;
    assign _16 = clock;
    assign _30 = _25 + _29;
    assign _27 = _25 == _26;
    assign _28 = ~ _27;
    assign _31 = _28 ? _30 : _25;
    assign _33 = _19 ? _32 : _31;
    assign _17 = _33;
    always @(posedge _16) begin
        _25 <= _17;
    end
    always @* begin
        case (_25)
        0: _90 <= _14;
        1: _90 <= _12;
        2: _90 <= _10;
        3: _90 <= _8;
        4: _90 <= _6;
        5: _90 <= _4;
        default: _90 <= _89;
        endcase
    end
    assign _19 = start_twiddles;
    assign _92 = _19 ? _91 : _90;
    assign _20 = _92;
    always @(posedge _16) begin
        _37 <= _20;
    end

    /* aliases */

    /* output assignments */
    assign w = _37;

endmodule
module dp (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_0 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1110000010010110111101100111110101000010010111011100100100000111;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0110111000001001111101011111101101111110101000111110001001000001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1001100001001110110001010001100101001101000000000101011100110101;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1001110110001111001010101101011110001011111111101101100101110010;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1001010001011000110101001011010000001101001101000000011100011110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0000011001010011101101001000000000011101101000011100100011001111;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1111001011000011010100011001100110010101100111011111110010110110;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_1 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1110111110011011001000010110000110000111101001101001011101000111;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0110000010000100111001101000010001011010100100010010111101001101;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0111101001011001000101011001010111100110011111000010011111101000;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0001100100000101110100000010101001011100010000010001111101001110;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0110111000001001111101011111101101111110101000111110001001000001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1001110110001111001010101101011110001011111111101101100101110010;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0000011001010011101101001000000000011101101000011100100011001111;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_2 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1110100111110010110110100110110010111110001000101100111000010001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0011101010100111000001000000100000001000111011011010110011010101;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1110000001000010100010111011011100101110110101110011010000101110;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0110000010000100111001101000010001011010100100010010111101001101;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1001110001100110000010001101010010111100110001111111101000100100;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0110111000001001111101011111101101111110101000111110001001000001;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1001010001011000110101001011010000001101001101000000011100011110;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_3 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0101010011010111101011100001010011111111011110000011001100001001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1011101000100101111010110101110011010001100101110000101011101011;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0011110110100000010111111110111001110000110001001111001010111010;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1011111101111001000101000011110011100110000011001010100101100110;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0110000010000100111001101000010001011010100100010010111101001101;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0001100100000101110100000010101001011100010000010001111101001110;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1001110110001111001010101101011110001011111111101101100101110010;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_4 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0111101110000001010101110000111011001001110000111111101100101101;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0000001101001101110010111010010110001010110001010000000000111110;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0100000000001010011100001110010111000101111110001100111000110011;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0011110110100000010111111110111001110000110001001111001010111010;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1110000001000010100010111011011100101110110101110011010000101110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0111101001011001000101011001010111100110011111000010011111101000;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1001100001001110110001010001100101001101000000000101011100110101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_5 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0110110110111110101101111110000000100110100001110010111000111001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1110010100001110110001011011010111010011000010010011010110000000;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0000001101001101110010111010010110001010110001010000000000111110;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1011101000100101111010110101110011010001100101110000101011101011;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0011101010100111000001000000100000001000111011011010110011010101;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0110000010000100111001101000010001011010100100010010111101001101;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0110111000001001111101011111101101111110101000111110001001000001;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_6 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1101011100010110100111110011100101110111000110010000001101000011;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0110110110111110101101111110000000100110100001110010111000111001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0111101110000001010101110000111011001001110000111111101100101101;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0101010011010111101011100001010011111111011110000011001100001001;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1110100111110010110110100110110010111110001000101100111000010001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1110111110011011001000010110000110000111101001101001011101000111;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1110000010010110111101100111110101000010010111011100100100000111;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module parallel_cores (
    wr_d7,
    wr_d6,
    wr_d5,
    wr_d4,
    wr_d3,
    wr_d2,
    wr_d1,
    wr_d0,
    wr_addr,
    wr_en,
    rd_addr,
    rd_en,
    flip,
    first_4step_pass,
    first_iter,
    start,
    clear,
    clock,
    done_,
    rd_q0,
    rd_q1,
    rd_q2,
    rd_q3,
    rd_q4,
    rd_q5,
    rd_q6,
    rd_q7
);

    input [63:0] wr_d7;
    input [63:0] wr_d6;
    input [63:0] wr_d5;
    input [63:0] wr_d4;
    input [63:0] wr_d3;
    input [63:0] wr_d2;
    input [63:0] wr_d1;
    input [63:0] wr_d0;
    input [5:0] wr_addr;
    input [7:0] wr_en;
    input [5:0] rd_addr;
    input [7:0] rd_en;
    input flip;
    input first_4step_pass;
    input first_iter;
    input start;
    input clear;
    input clock;
    output done_;
    output [63:0] rd_q0;
    output [63:0] rd_q1;
    output [63:0] rd_q2;
    output [63:0] rd_q3;
    output [63:0] rd_q4;
    output [63:0] rd_q5;
    output [63:0] rd_q6;
    output [63:0] rd_q7;

    /* signal declarations */
    wire [5:0] address;
    wire write_enable;
    wire [5:0] address_0;
    wire _362;
    wire read_enable;
    wire _360;
    wire write_enable_0;
    wire _364;
    wire [131:0] _369;
    wire [63:0] _370;
    wire [5:0] _355 = 6'b000000;
    wire [5:0] address_1;
    wire _353;
    wire write_enable_1;
    wire [63:0] _267;
    wire [63:0] _266;
    wire [63:0] _268;
    wire [63:0] _264;
    wire [63:0] _263;
    wire [63:0] q1;
    wire [63:0] _269;
    wire [5:0] address_2;
    wire write_enable_2 = 1'b0;
    wire _254;
    wire read_enable_0;
    wire [5:0] address_3;
    wire _250;
    wire read_enable_1;
    wire _248;
    wire write_enable_3;
    wire _252;
    wire [131:0] _259;
    wire [63:0] _260;
    wire [63:0] data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_0;
    wire [5:0] _242 = 6'b000000;
    wire _240;
    wire _239;
    wire _238;
    wire _237;
    wire _236;
    wire _235;
    wire [5:0] _241;
    wire [5:0] address_4;
    wire write_enable_4 = 1'b0;
    wire _232;
    wire read_enable_2;
    wire [63:0] data_1;
    wire [63:0] data_2;
    wire _229;
    wire _228;
    wire _227;
    wire _226;
    wire _225;
    wire _224;
    wire [5:0] _230;
    wire [5:0] address_5;
    wire _221;
    wire read_enable_3;
    wire _219;
    wire write_enable_5;
    wire _223;
    wire [131:0] _246;
    wire [63:0] _247;
    wire _87 = 1'b0;
    wire _86 = 1'b0;
    wire _89;
    wire _3;
    reg PHASE;
    wire [63:0] _261;
    wire [5:0] address_6;
    wire _211;
    wire read_enable_4;
    wire write_enable_6;
    wire _213;
    wire [5:0] address_7;
    wire _206;
    wire read_enable_5;
    wire _204;
    wire write_enable_7;
    wire _208;
    wire [131:0] _216;
    wire [63:0] _217;
    wire [63:0] _283;
    wire [63:0] data_3;
    wire [63:0] data_4;
    wire [63:0] data_5;
    wire [63:0] data_6;
    wire [5:0] address_8;
    wire _169;
    wire read_enable_6;
    wire _166;
    wire _167;
    wire write_enable_8;
    wire _171;
    wire [5:0] address_9;
    wire _134;
    wire read_enable_7;
    wire _131;
    wire _132;
    wire write_enable_9;
    wire _136;
    wire [131:0] _202;
    wire [63:0] _203;
    wire _98 = 1'b0;
    wire _97 = 1'b0;
    wire _284;
    wire _5;
    reg PHASE_0;
    wire [63:0] q0;
    wire _94 = 1'b0;
    wire _93 = 1'b0;
    reg _96;
    wire [63:0] _262;
    wire [191:0] _282;
    wire [63:0] _285;
    wire [63:0] data_7;
    wire [63:0] data_8;
    wire [63:0] data_9;
    wire [63:0] data_10;
    wire [5:0] address_10;
    wire _349;
    wire _348;
    wire read_enable_8;
    wire _342 = 1'b0;
    wire _341 = 1'b0;
    wire _339 = 1'b0;
    wire _338 = 1'b0;
    wire _336 = 1'b0;
    wire _335 = 1'b0;
    wire _333 = 1'b0;
    wire _332 = 1'b0;
    wire _330 = 1'b0;
    wire _329 = 1'b0;
    wire _327 = 1'b0;
    wire _326 = 1'b0;
    wire _324 = 1'b0;
    wire _323 = 1'b0;
    wire _321 = 1'b0;
    wire _320 = 1'b0;
    wire _318 = 1'b0;
    wire _317 = 1'b0;
    reg _319;
    reg _322;
    reg _325;
    reg _328;
    reg _331;
    reg _334;
    reg _337;
    reg _340;
    reg _343;
    wire _344;
    wire _315 = 1'b0;
    wire _314 = 1'b0;
    wire _312 = 1'b0;
    wire _311 = 1'b0;
    wire _309 = 1'b0;
    wire _308 = 1'b0;
    wire _306 = 1'b0;
    wire _305 = 1'b0;
    wire _303 = 1'b0;
    wire _302 = 1'b0;
    wire _300 = 1'b0;
    wire _299 = 1'b0;
    wire _297 = 1'b0;
    wire _296 = 1'b0;
    wire _294 = 1'b0;
    wire _293 = 1'b0;
    wire _291 = 1'b0;
    wire _290 = 1'b0;
    reg _292;
    reg _295;
    reg _298;
    reg _301;
    reg _304;
    reg _307;
    reg _310;
    reg _313;
    reg _316;
    wire _345;
    wire _346;
    wire write_enable_10;
    wire _351;
    wire [131:0] _358;
    wire [63:0] _359;
    wire _287 = 1'b0;
    wire _286 = 1'b0;
    wire _289;
    wire _7;
    reg PHASE_1;
    wire [63:0] _371;
    wire [5:0] address_11;
    wire write_enable_11;
    wire [5:0] address_12;
    wire _546;
    wire read_enable_9;
    wire _544;
    wire write_enable_12;
    wire _548;
    wire [131:0] _553;
    wire [63:0] _554;
    wire [5:0] _539 = 6'b000000;
    wire [5:0] address_13;
    wire _537;
    wire write_enable_13;
    wire [63:0] _462;
    wire [63:0] _461;
    wire [63:0] _463;
    wire [63:0] _459;
    wire [63:0] _458;
    wire [63:0] q1_0;
    wire [63:0] _464;
    wire [5:0] address_14;
    wire write_enable_14 = 1'b0;
    wire _449;
    wire read_enable_10;
    wire [5:0] address_15;
    wire _445;
    wire read_enable_11;
    wire _443;
    wire write_enable_15;
    wire _447;
    wire [131:0] _454;
    wire [63:0] _455;
    wire [63:0] data_11 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_12;
    wire [5:0] _437 = 6'b000000;
    wire _435;
    wire _434;
    wire _433;
    wire _432;
    wire _431;
    wire _430;
    wire [5:0] _436;
    wire [5:0] address_16;
    wire write_enable_16 = 1'b0;
    wire _427;
    wire read_enable_12;
    wire [63:0] data_13;
    wire [63:0] data_14;
    wire _424;
    wire _423;
    wire _422;
    wire _421;
    wire _420;
    wire _419;
    wire [5:0] _425;
    wire [5:0] address_17;
    wire _416;
    wire read_enable_13;
    wire _414;
    wire write_enable_17;
    wire _418;
    wire [131:0] _441;
    wire [63:0] _442;
    wire _373 = 1'b0;
    wire _372 = 1'b0;
    wire _375;
    wire _11;
    reg PHASE_2;
    wire [63:0] _456;
    wire [5:0] address_18;
    wire _406;
    wire read_enable_14;
    wire write_enable_18;
    wire _408;
    wire [5:0] address_19;
    wire _401;
    wire read_enable_15;
    wire _399;
    wire write_enable_19;
    wire _403;
    wire [131:0] _411;
    wire [63:0] _412;
    wire [63:0] _467;
    wire [63:0] data_15;
    wire [63:0] data_16;
    wire [63:0] data_17;
    wire [63:0] data_18;
    wire [5:0] address_20;
    wire _392;
    wire read_enable_16;
    wire _389;
    wire _390;
    wire write_enable_20;
    wire _394;
    wire [5:0] address_21;
    wire _385;
    wire read_enable_17;
    wire _382;
    wire _383;
    wire write_enable_21;
    wire _387;
    wire [131:0] _397;
    wire [63:0] _398;
    wire _380 = 1'b0;
    wire _379 = 1'b0;
    wire _468;
    wire _13;
    reg PHASE_3;
    wire [63:0] q0_0;
    wire _377 = 1'b0;
    wire _376 = 1'b0;
    reg _378;
    wire [63:0] _457;
    wire [191:0] _466;
    wire [63:0] _469;
    wire [63:0] data_19;
    wire [63:0] data_20;
    wire [63:0] data_21;
    wire [63:0] data_22;
    wire [5:0] address_22;
    wire _533;
    wire _532;
    wire read_enable_18;
    wire _526 = 1'b0;
    wire _525 = 1'b0;
    wire _523 = 1'b0;
    wire _522 = 1'b0;
    wire _520 = 1'b0;
    wire _519 = 1'b0;
    wire _517 = 1'b0;
    wire _516 = 1'b0;
    wire _514 = 1'b0;
    wire _513 = 1'b0;
    wire _511 = 1'b0;
    wire _510 = 1'b0;
    wire _508 = 1'b0;
    wire _507 = 1'b0;
    wire _505 = 1'b0;
    wire _504 = 1'b0;
    wire _502 = 1'b0;
    wire _501 = 1'b0;
    reg _503;
    reg _506;
    reg _509;
    reg _512;
    reg _515;
    reg _518;
    reg _521;
    reg _524;
    reg _527;
    wire _528;
    wire _499 = 1'b0;
    wire _498 = 1'b0;
    wire _496 = 1'b0;
    wire _495 = 1'b0;
    wire _493 = 1'b0;
    wire _492 = 1'b0;
    wire _490 = 1'b0;
    wire _489 = 1'b0;
    wire _487 = 1'b0;
    wire _486 = 1'b0;
    wire _484 = 1'b0;
    wire _483 = 1'b0;
    wire _481 = 1'b0;
    wire _480 = 1'b0;
    wire _478 = 1'b0;
    wire _477 = 1'b0;
    wire _475 = 1'b0;
    wire _474 = 1'b0;
    reg _476;
    reg _479;
    reg _482;
    reg _485;
    reg _488;
    reg _491;
    reg _494;
    reg _497;
    reg _500;
    wire _529;
    wire _530;
    wire write_enable_22;
    wire _535;
    wire [131:0] _542;
    wire [63:0] _543;
    wire _471 = 1'b0;
    wire _470 = 1'b0;
    wire _473;
    wire _15;
    reg PHASE_4;
    wire [63:0] _555;
    wire [5:0] address_23;
    wire write_enable_23;
    wire [5:0] address_24;
    wire _730;
    wire read_enable_19;
    wire _728;
    wire write_enable_24;
    wire _732;
    wire [131:0] _737;
    wire [63:0] _738;
    wire [5:0] _723 = 6'b000000;
    wire [5:0] address_25;
    wire _721;
    wire write_enable_25;
    wire [63:0] _646;
    wire [63:0] _645;
    wire [63:0] _647;
    wire [63:0] _643;
    wire [63:0] _642;
    wire [63:0] q1_1;
    wire [63:0] _648;
    wire [5:0] address_26;
    wire write_enable_26 = 1'b0;
    wire _633;
    wire read_enable_20;
    wire [5:0] address_27;
    wire _629;
    wire read_enable_21;
    wire _627;
    wire write_enable_27;
    wire _631;
    wire [131:0] _638;
    wire [63:0] _639;
    wire [63:0] data_23 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_24;
    wire [5:0] _621 = 6'b000000;
    wire _619;
    wire _618;
    wire _617;
    wire _616;
    wire _615;
    wire _614;
    wire [5:0] _620;
    wire [5:0] address_28;
    wire write_enable_28 = 1'b0;
    wire _611;
    wire read_enable_22;
    wire [63:0] data_25;
    wire [63:0] data_26;
    wire _608;
    wire _607;
    wire _606;
    wire _605;
    wire _604;
    wire _603;
    wire [5:0] _609;
    wire [5:0] address_29;
    wire _600;
    wire read_enable_23;
    wire _598;
    wire write_enable_29;
    wire _602;
    wire [131:0] _625;
    wire [63:0] _626;
    wire _557 = 1'b0;
    wire _556 = 1'b0;
    wire _559;
    wire _19;
    reg PHASE_5;
    wire [63:0] _640;
    wire [5:0] address_30;
    wire _590;
    wire read_enable_24;
    wire write_enable_30;
    wire _592;
    wire [5:0] address_31;
    wire _585;
    wire read_enable_25;
    wire _583;
    wire write_enable_31;
    wire _587;
    wire [131:0] _595;
    wire [63:0] _596;
    wire [63:0] _651;
    wire [63:0] data_27;
    wire [63:0] data_28;
    wire [63:0] data_29;
    wire [63:0] data_30;
    wire [5:0] address_32;
    wire _576;
    wire read_enable_26;
    wire _573;
    wire _574;
    wire write_enable_32;
    wire _578;
    wire [5:0] address_33;
    wire _569;
    wire read_enable_27;
    wire _566;
    wire _567;
    wire write_enable_33;
    wire _571;
    wire [131:0] _581;
    wire [63:0] _582;
    wire _564 = 1'b0;
    wire _563 = 1'b0;
    wire _652;
    wire _21;
    reg PHASE_6;
    wire [63:0] q0_1;
    wire _561 = 1'b0;
    wire _560 = 1'b0;
    reg _562;
    wire [63:0] _641;
    wire [191:0] _650;
    wire [63:0] _653;
    wire [63:0] data_31;
    wire [63:0] data_32;
    wire [63:0] data_33;
    wire [63:0] data_34;
    wire [5:0] address_34;
    wire _717;
    wire _716;
    wire read_enable_28;
    wire _710 = 1'b0;
    wire _709 = 1'b0;
    wire _707 = 1'b0;
    wire _706 = 1'b0;
    wire _704 = 1'b0;
    wire _703 = 1'b0;
    wire _701 = 1'b0;
    wire _700 = 1'b0;
    wire _698 = 1'b0;
    wire _697 = 1'b0;
    wire _695 = 1'b0;
    wire _694 = 1'b0;
    wire _692 = 1'b0;
    wire _691 = 1'b0;
    wire _689 = 1'b0;
    wire _688 = 1'b0;
    wire _686 = 1'b0;
    wire _685 = 1'b0;
    reg _687;
    reg _690;
    reg _693;
    reg _696;
    reg _699;
    reg _702;
    reg _705;
    reg _708;
    reg _711;
    wire _712;
    wire _683 = 1'b0;
    wire _682 = 1'b0;
    wire _680 = 1'b0;
    wire _679 = 1'b0;
    wire _677 = 1'b0;
    wire _676 = 1'b0;
    wire _674 = 1'b0;
    wire _673 = 1'b0;
    wire _671 = 1'b0;
    wire _670 = 1'b0;
    wire _668 = 1'b0;
    wire _667 = 1'b0;
    wire _665 = 1'b0;
    wire _664 = 1'b0;
    wire _662 = 1'b0;
    wire _661 = 1'b0;
    wire _659 = 1'b0;
    wire _658 = 1'b0;
    reg _660;
    reg _663;
    reg _666;
    reg _669;
    reg _672;
    reg _675;
    reg _678;
    reg _681;
    reg _684;
    wire _713;
    wire _714;
    wire write_enable_34;
    wire _719;
    wire [131:0] _726;
    wire [63:0] _727;
    wire _655 = 1'b0;
    wire _654 = 1'b0;
    wire _657;
    wire _23;
    reg PHASE_7;
    wire [63:0] _739;
    wire [5:0] address_35;
    wire write_enable_35;
    wire [5:0] address_36;
    wire _914;
    wire read_enable_29;
    wire _912;
    wire write_enable_36;
    wire _916;
    wire [131:0] _921;
    wire [63:0] _922;
    wire [5:0] _907 = 6'b000000;
    wire [5:0] address_37;
    wire _905;
    wire write_enable_37;
    wire [63:0] _830;
    wire [63:0] _829;
    wire [63:0] _831;
    wire [63:0] _827;
    wire [63:0] _826;
    wire [63:0] q1_2;
    wire [63:0] _832;
    wire [5:0] address_38;
    wire write_enable_38 = 1'b0;
    wire _817;
    wire read_enable_30;
    wire [5:0] address_39;
    wire _813;
    wire read_enable_31;
    wire _811;
    wire write_enable_39;
    wire _815;
    wire [131:0] _822;
    wire [63:0] _823;
    wire [63:0] data_35 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_36;
    wire [5:0] _805 = 6'b000000;
    wire _803;
    wire _802;
    wire _801;
    wire _800;
    wire _799;
    wire _798;
    wire [5:0] _804;
    wire [5:0] address_40;
    wire write_enable_40 = 1'b0;
    wire _795;
    wire read_enable_32;
    wire [63:0] data_37;
    wire [63:0] data_38;
    wire _792;
    wire _791;
    wire _790;
    wire _789;
    wire _788;
    wire _787;
    wire [5:0] _793;
    wire [5:0] address_41;
    wire _784;
    wire read_enable_33;
    wire _782;
    wire write_enable_41;
    wire _786;
    wire [131:0] _809;
    wire [63:0] _810;
    wire _741 = 1'b0;
    wire _740 = 1'b0;
    wire _743;
    wire _27;
    reg PHASE_8;
    wire [63:0] _824;
    wire [5:0] address_42;
    wire _774;
    wire read_enable_34;
    wire write_enable_42;
    wire _776;
    wire [5:0] address_43;
    wire _769;
    wire read_enable_35;
    wire _767;
    wire write_enable_43;
    wire _771;
    wire [131:0] _779;
    wire [63:0] _780;
    wire [63:0] _835;
    wire [63:0] data_39;
    wire [63:0] data_40;
    wire [63:0] data_41;
    wire [63:0] data_42;
    wire [5:0] address_44;
    wire _760;
    wire read_enable_36;
    wire _757;
    wire _758;
    wire write_enable_44;
    wire _762;
    wire [5:0] address_45;
    wire _753;
    wire read_enable_37;
    wire _750;
    wire _751;
    wire write_enable_45;
    wire _755;
    wire [131:0] _765;
    wire [63:0] _766;
    wire _748 = 1'b0;
    wire _747 = 1'b0;
    wire _836;
    wire _29;
    reg PHASE_9;
    wire [63:0] q0_2;
    wire _745 = 1'b0;
    wire _744 = 1'b0;
    reg _746;
    wire [63:0] _825;
    wire [191:0] _834;
    wire [63:0] _837;
    wire [63:0] data_43;
    wire [63:0] data_44;
    wire [63:0] data_45;
    wire [63:0] data_46;
    wire [5:0] address_46;
    wire _901;
    wire _900;
    wire read_enable_38;
    wire _894 = 1'b0;
    wire _893 = 1'b0;
    wire _891 = 1'b0;
    wire _890 = 1'b0;
    wire _888 = 1'b0;
    wire _887 = 1'b0;
    wire _885 = 1'b0;
    wire _884 = 1'b0;
    wire _882 = 1'b0;
    wire _881 = 1'b0;
    wire _879 = 1'b0;
    wire _878 = 1'b0;
    wire _876 = 1'b0;
    wire _875 = 1'b0;
    wire _873 = 1'b0;
    wire _872 = 1'b0;
    wire _870 = 1'b0;
    wire _869 = 1'b0;
    reg _871;
    reg _874;
    reg _877;
    reg _880;
    reg _883;
    reg _886;
    reg _889;
    reg _892;
    reg _895;
    wire _896;
    wire _867 = 1'b0;
    wire _866 = 1'b0;
    wire _864 = 1'b0;
    wire _863 = 1'b0;
    wire _861 = 1'b0;
    wire _860 = 1'b0;
    wire _858 = 1'b0;
    wire _857 = 1'b0;
    wire _855 = 1'b0;
    wire _854 = 1'b0;
    wire _852 = 1'b0;
    wire _851 = 1'b0;
    wire _849 = 1'b0;
    wire _848 = 1'b0;
    wire _846 = 1'b0;
    wire _845 = 1'b0;
    wire _843 = 1'b0;
    wire _842 = 1'b0;
    reg _844;
    reg _847;
    reg _850;
    reg _853;
    reg _856;
    reg _859;
    reg _862;
    reg _865;
    reg _868;
    wire _897;
    wire _898;
    wire write_enable_46;
    wire _903;
    wire [131:0] _910;
    wire [63:0] _911;
    wire _839 = 1'b0;
    wire _838 = 1'b0;
    wire _841;
    wire _31;
    reg PHASE_10;
    wire [63:0] _923;
    wire [5:0] address_47;
    wire write_enable_47;
    wire [5:0] address_48;
    wire _1098;
    wire read_enable_39;
    wire _1096;
    wire write_enable_48;
    wire _1100;
    wire [131:0] _1105;
    wire [63:0] _1106;
    wire [5:0] _1091 = 6'b000000;
    wire [5:0] address_49;
    wire _1089;
    wire write_enable_49;
    wire [63:0] _1014;
    wire [63:0] _1013;
    wire [63:0] _1015;
    wire [63:0] _1011;
    wire [63:0] _1010;
    wire [63:0] q1_3;
    wire [63:0] _1016;
    wire [5:0] address_50;
    wire write_enable_50 = 1'b0;
    wire _1001;
    wire read_enable_40;
    wire [5:0] address_51;
    wire _997;
    wire read_enable_41;
    wire _995;
    wire write_enable_51;
    wire _999;
    wire [131:0] _1006;
    wire [63:0] _1007;
    wire [63:0] data_47 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_48;
    wire [5:0] _989 = 6'b000000;
    wire _987;
    wire _986;
    wire _985;
    wire _984;
    wire _983;
    wire _982;
    wire [5:0] _988;
    wire [5:0] address_52;
    wire write_enable_52 = 1'b0;
    wire _979;
    wire read_enable_42;
    wire [63:0] data_49;
    wire [63:0] data_50;
    wire _976;
    wire _975;
    wire _974;
    wire _973;
    wire _972;
    wire _971;
    wire [5:0] _977;
    wire [5:0] address_53;
    wire _968;
    wire read_enable_43;
    wire _966;
    wire write_enable_53;
    wire _970;
    wire [131:0] _993;
    wire [63:0] _994;
    wire _925 = 1'b0;
    wire _924 = 1'b0;
    wire _927;
    wire _35;
    reg PHASE_11;
    wire [63:0] _1008;
    wire [5:0] address_54;
    wire _958;
    wire read_enable_44;
    wire write_enable_54;
    wire _960;
    wire [5:0] address_55;
    wire _953;
    wire read_enable_45;
    wire _951;
    wire write_enable_55;
    wire _955;
    wire [131:0] _963;
    wire [63:0] _964;
    wire [63:0] _1019;
    wire [63:0] data_51;
    wire [63:0] data_52;
    wire [63:0] data_53;
    wire [63:0] data_54;
    wire [5:0] address_56;
    wire _944;
    wire read_enable_46;
    wire _941;
    wire _942;
    wire write_enable_56;
    wire _946;
    wire [5:0] address_57;
    wire _937;
    wire read_enable_47;
    wire _934;
    wire _935;
    wire write_enable_57;
    wire _939;
    wire [131:0] _949;
    wire [63:0] _950;
    wire _932 = 1'b0;
    wire _931 = 1'b0;
    wire _1020;
    wire _37;
    reg PHASE_12;
    wire [63:0] q0_3;
    wire _929 = 1'b0;
    wire _928 = 1'b0;
    reg _930;
    wire [63:0] _1009;
    wire [191:0] _1018;
    wire [63:0] _1021;
    wire [63:0] data_55;
    wire [63:0] data_56;
    wire [63:0] data_57;
    wire [63:0] data_58;
    wire [5:0] address_58;
    wire _1085;
    wire _1084;
    wire read_enable_48;
    wire _1078 = 1'b0;
    wire _1077 = 1'b0;
    wire _1075 = 1'b0;
    wire _1074 = 1'b0;
    wire _1072 = 1'b0;
    wire _1071 = 1'b0;
    wire _1069 = 1'b0;
    wire _1068 = 1'b0;
    wire _1066 = 1'b0;
    wire _1065 = 1'b0;
    wire _1063 = 1'b0;
    wire _1062 = 1'b0;
    wire _1060 = 1'b0;
    wire _1059 = 1'b0;
    wire _1057 = 1'b0;
    wire _1056 = 1'b0;
    wire _1054 = 1'b0;
    wire _1053 = 1'b0;
    reg _1055;
    reg _1058;
    reg _1061;
    reg _1064;
    reg _1067;
    reg _1070;
    reg _1073;
    reg _1076;
    reg _1079;
    wire _1080;
    wire _1051 = 1'b0;
    wire _1050 = 1'b0;
    wire _1048 = 1'b0;
    wire _1047 = 1'b0;
    wire _1045 = 1'b0;
    wire _1044 = 1'b0;
    wire _1042 = 1'b0;
    wire _1041 = 1'b0;
    wire _1039 = 1'b0;
    wire _1038 = 1'b0;
    wire _1036 = 1'b0;
    wire _1035 = 1'b0;
    wire _1033 = 1'b0;
    wire _1032 = 1'b0;
    wire _1030 = 1'b0;
    wire _1029 = 1'b0;
    wire _1027 = 1'b0;
    wire _1026 = 1'b0;
    reg _1028;
    reg _1031;
    reg _1034;
    reg _1037;
    reg _1040;
    reg _1043;
    reg _1046;
    reg _1049;
    reg _1052;
    wire _1081;
    wire _1082;
    wire write_enable_58;
    wire _1087;
    wire [131:0] _1094;
    wire [63:0] _1095;
    wire _1023 = 1'b0;
    wire _1022 = 1'b0;
    wire _1025;
    wire _39;
    reg PHASE_13;
    wire [63:0] _1107;
    wire [5:0] address_59;
    wire write_enable_59;
    wire [5:0] address_60;
    wire _1282;
    wire read_enable_49;
    wire _1280;
    wire write_enable_60;
    wire _1284;
    wire [131:0] _1289;
    wire [63:0] _1290;
    wire [5:0] _1275 = 6'b000000;
    wire [5:0] address_61;
    wire _1273;
    wire write_enable_61;
    wire [63:0] _1198;
    wire [63:0] _1197;
    wire [63:0] _1199;
    wire [63:0] _1195;
    wire [63:0] _1194;
    wire [63:0] q1_4;
    wire [63:0] _1200;
    wire [5:0] address_62;
    wire write_enable_62 = 1'b0;
    wire _1185;
    wire read_enable_50;
    wire [5:0] address_63;
    wire _1181;
    wire read_enable_51;
    wire _1179;
    wire write_enable_63;
    wire _1183;
    wire [131:0] _1190;
    wire [63:0] _1191;
    wire [63:0] data_59 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_60;
    wire [5:0] _1173 = 6'b000000;
    wire _1171;
    wire _1170;
    wire _1169;
    wire _1168;
    wire _1167;
    wire _1166;
    wire [5:0] _1172;
    wire [5:0] address_64;
    wire write_enable_64 = 1'b0;
    wire _1163;
    wire read_enable_52;
    wire [63:0] data_61;
    wire [63:0] data_62;
    wire _1160;
    wire _1159;
    wire _1158;
    wire _1157;
    wire _1156;
    wire _1155;
    wire [5:0] _1161;
    wire [5:0] address_65;
    wire _1152;
    wire read_enable_53;
    wire _1150;
    wire write_enable_65;
    wire _1154;
    wire [131:0] _1177;
    wire [63:0] _1178;
    wire _1109 = 1'b0;
    wire _1108 = 1'b0;
    wire _1111;
    wire _43;
    reg PHASE_14;
    wire [63:0] _1192;
    wire [5:0] address_66;
    wire _1142;
    wire read_enable_54;
    wire write_enable_66;
    wire _1144;
    wire [5:0] address_67;
    wire _1137;
    wire read_enable_55;
    wire _1135;
    wire write_enable_67;
    wire _1139;
    wire [131:0] _1147;
    wire [63:0] _1148;
    wire [63:0] _1203;
    wire [63:0] data_63;
    wire [63:0] data_64;
    wire [63:0] data_65;
    wire [63:0] data_66;
    wire [5:0] address_68;
    wire _1128;
    wire read_enable_56;
    wire _1125;
    wire _1126;
    wire write_enable_68;
    wire _1130;
    wire [5:0] address_69;
    wire _1121;
    wire read_enable_57;
    wire _1118;
    wire _1119;
    wire write_enable_69;
    wire _1123;
    wire [131:0] _1133;
    wire [63:0] _1134;
    wire _1116 = 1'b0;
    wire _1115 = 1'b0;
    wire _1204;
    wire _45;
    reg PHASE_15;
    wire [63:0] q0_4;
    wire _1113 = 1'b0;
    wire _1112 = 1'b0;
    reg _1114;
    wire [63:0] _1193;
    wire [191:0] _1202;
    wire [63:0] _1205;
    wire [63:0] data_67;
    wire [63:0] data_68;
    wire [63:0] data_69;
    wire [63:0] data_70;
    wire [5:0] address_70;
    wire _1269;
    wire _1268;
    wire read_enable_58;
    wire _1262 = 1'b0;
    wire _1261 = 1'b0;
    wire _1259 = 1'b0;
    wire _1258 = 1'b0;
    wire _1256 = 1'b0;
    wire _1255 = 1'b0;
    wire _1253 = 1'b0;
    wire _1252 = 1'b0;
    wire _1250 = 1'b0;
    wire _1249 = 1'b0;
    wire _1247 = 1'b0;
    wire _1246 = 1'b0;
    wire _1244 = 1'b0;
    wire _1243 = 1'b0;
    wire _1241 = 1'b0;
    wire _1240 = 1'b0;
    wire _1238 = 1'b0;
    wire _1237 = 1'b0;
    reg _1239;
    reg _1242;
    reg _1245;
    reg _1248;
    reg _1251;
    reg _1254;
    reg _1257;
    reg _1260;
    reg _1263;
    wire _1264;
    wire _1235 = 1'b0;
    wire _1234 = 1'b0;
    wire _1232 = 1'b0;
    wire _1231 = 1'b0;
    wire _1229 = 1'b0;
    wire _1228 = 1'b0;
    wire _1226 = 1'b0;
    wire _1225 = 1'b0;
    wire _1223 = 1'b0;
    wire _1222 = 1'b0;
    wire _1220 = 1'b0;
    wire _1219 = 1'b0;
    wire _1217 = 1'b0;
    wire _1216 = 1'b0;
    wire _1214 = 1'b0;
    wire _1213 = 1'b0;
    wire _1211 = 1'b0;
    wire _1210 = 1'b0;
    reg _1212;
    reg _1215;
    reg _1218;
    reg _1221;
    reg _1224;
    reg _1227;
    reg _1230;
    reg _1233;
    reg _1236;
    wire _1265;
    wire _1266;
    wire write_enable_70;
    wire _1271;
    wire [131:0] _1278;
    wire [63:0] _1279;
    wire _1207 = 1'b0;
    wire _1206 = 1'b0;
    wire _1209;
    wire _47;
    reg PHASE_16;
    wire [63:0] _1291;
    wire [5:0] address_71;
    wire write_enable_71;
    wire [5:0] address_72;
    wire _1466;
    wire read_enable_59;
    wire _1464;
    wire write_enable_72;
    wire _1468;
    wire [131:0] _1473;
    wire [63:0] _1474;
    wire [5:0] _1459 = 6'b000000;
    wire [5:0] address_73;
    wire _1457;
    wire write_enable_73;
    wire [63:0] _1382;
    wire [63:0] _1381;
    wire [63:0] _1383;
    wire [63:0] _1379;
    wire [63:0] _1378;
    wire [63:0] q1_5;
    wire [63:0] _1384;
    wire [5:0] address_74;
    wire write_enable_74 = 1'b0;
    wire _1369;
    wire read_enable_60;
    wire [5:0] address_75;
    wire _1365;
    wire read_enable_61;
    wire _1363;
    wire write_enable_75;
    wire _1367;
    wire [131:0] _1374;
    wire [63:0] _1375;
    wire [63:0] data_71 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_72;
    wire [5:0] _1357 = 6'b000000;
    wire _1355;
    wire _1354;
    wire _1353;
    wire _1352;
    wire _1351;
    wire _1350;
    wire [5:0] _1356;
    wire [5:0] address_76;
    wire write_enable_76 = 1'b0;
    wire _1347;
    wire read_enable_62;
    wire [63:0] data_73;
    wire [63:0] data_74;
    wire _1344;
    wire _1343;
    wire _1342;
    wire _1341;
    wire _1340;
    wire _1339;
    wire [5:0] _1345;
    wire [5:0] address_77;
    wire _1336;
    wire read_enable_63;
    wire _1334;
    wire write_enable_77;
    wire _1338;
    wire [131:0] _1361;
    wire [63:0] _1362;
    wire _1293 = 1'b0;
    wire _1292 = 1'b0;
    wire _1295;
    wire _51;
    reg PHASE_17;
    wire [63:0] _1376;
    wire [5:0] address_78;
    wire _1326;
    wire read_enable_64;
    wire write_enable_78;
    wire _1328;
    wire [5:0] address_79;
    wire _1321;
    wire read_enable_65;
    wire _1319;
    wire write_enable_79;
    wire _1323;
    wire [131:0] _1331;
    wire [63:0] _1332;
    wire [63:0] _1387;
    wire [63:0] data_75;
    wire [63:0] data_76;
    wire [63:0] data_77;
    wire [63:0] data_78;
    wire [5:0] address_80;
    wire _1312;
    wire read_enable_66;
    wire _1309;
    wire _1310;
    wire write_enable_80;
    wire _1314;
    wire [5:0] address_81;
    wire _1305;
    wire read_enable_67;
    wire _1302;
    wire _1303;
    wire write_enable_81;
    wire _1307;
    wire [131:0] _1317;
    wire [63:0] _1318;
    wire _1300 = 1'b0;
    wire _1299 = 1'b0;
    wire _1388;
    wire _53;
    reg PHASE_18;
    wire [63:0] q0_5;
    wire _1297 = 1'b0;
    wire _1296 = 1'b0;
    reg _1298;
    wire [63:0] _1377;
    wire [191:0] _1386;
    wire [63:0] _1389;
    wire [63:0] data_79;
    wire [63:0] data_80;
    wire [63:0] data_81;
    wire [63:0] data_82;
    wire [5:0] address_82;
    wire _1453;
    wire _1452;
    wire read_enable_68;
    wire _1446 = 1'b0;
    wire _1445 = 1'b0;
    wire _1443 = 1'b0;
    wire _1442 = 1'b0;
    wire _1440 = 1'b0;
    wire _1439 = 1'b0;
    wire _1437 = 1'b0;
    wire _1436 = 1'b0;
    wire _1434 = 1'b0;
    wire _1433 = 1'b0;
    wire _1431 = 1'b0;
    wire _1430 = 1'b0;
    wire _1428 = 1'b0;
    wire _1427 = 1'b0;
    wire _1425 = 1'b0;
    wire _1424 = 1'b0;
    wire _1422 = 1'b0;
    wire _1421 = 1'b0;
    reg _1423;
    reg _1426;
    reg _1429;
    reg _1432;
    reg _1435;
    reg _1438;
    reg _1441;
    reg _1444;
    reg _1447;
    wire _1448;
    wire _1419 = 1'b0;
    wire _1418 = 1'b0;
    wire _1416 = 1'b0;
    wire _1415 = 1'b0;
    wire _1413 = 1'b0;
    wire _1412 = 1'b0;
    wire _1410 = 1'b0;
    wire _1409 = 1'b0;
    wire _1407 = 1'b0;
    wire _1406 = 1'b0;
    wire _1404 = 1'b0;
    wire _1403 = 1'b0;
    wire _1401 = 1'b0;
    wire _1400 = 1'b0;
    wire _1398 = 1'b0;
    wire _1397 = 1'b0;
    wire _1395 = 1'b0;
    wire _1394 = 1'b0;
    reg _1396;
    reg _1399;
    reg _1402;
    reg _1405;
    reg _1408;
    reg _1411;
    reg _1414;
    reg _1417;
    reg _1420;
    wire _1449;
    wire _1450;
    wire write_enable_82;
    wire _1455;
    wire [131:0] _1462;
    wire [63:0] _1463;
    wire _1391 = 1'b0;
    wire _1390 = 1'b0;
    wire _1393;
    wire _55;
    reg PHASE_19;
    wire [63:0] _1475;
    wire [5:0] address_83;
    wire write_enable_83;
    wire [5:0] address_84;
    wire _1650;
    wire read_enable_69;
    wire _1648;
    wire write_enable_84;
    wire _1652;
    wire [131:0] _1657;
    wire [63:0] _1658;
    wire [5:0] _1643 = 6'b000000;
    wire [5:0] address_85;
    wire _1641;
    wire write_enable_85;
    wire [3:0] _280;
    wire _279;
    wire _277;
    wire [63:0] _276;
    wire [63:0] _275;
    wire [63:0] _274;
    wire [63:0] _273;
    wire [63:0] _272;
    wire [63:0] _271;
    wire [63:0] _270;
    wire [63:0] _1566;
    wire [63:0] _1565;
    wire [63:0] _1567;
    wire [63:0] _1563;
    wire [63:0] _1562;
    wire [63:0] q1_6;
    wire [63:0] _1568;
    wire [5:0] address_86;
    wire write_enable_86 = 1'b0;
    wire _1553;
    wire read_enable_70;
    wire [5:0] address_87;
    wire _1549;
    wire read_enable_71;
    wire _1547;
    wire write_enable_87;
    wire _1551;
    wire [131:0] _1558;
    wire [63:0] _1559;
    wire [63:0] data_83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_84;
    wire [5:0] _1541 = 6'b000000;
    wire _1539;
    wire _1538;
    wire _1537;
    wire _1536;
    wire _1535;
    wire _1534;
    wire [5:0] _1540;
    wire [5:0] address_88;
    wire write_enable_88 = 1'b0;
    wire _1531;
    wire read_enable_72;
    wire [63:0] data_85;
    wire [63:0] data_86;
    wire [5:0] _60;
    wire _1528;
    wire _1527;
    wire _1526;
    wire _1525;
    wire _1524;
    wire _1523;
    wire [5:0] _1529;
    wire [5:0] address_89;
    wire _1520;
    wire read_enable_73;
    wire [7:0] _62;
    wire _1518;
    wire write_enable_89;
    wire _1522;
    wire [131:0] _1545;
    wire [63:0] _1546;
    wire _1477 = 1'b0;
    wire _1476 = 1'b0;
    wire _1479;
    wire _63;
    reg PHASE_20;
    wire [63:0] _1560;
    wire [5:0] address_90;
    wire _1510;
    wire read_enable_74;
    wire write_enable_90;
    wire _1512;
    wire [5:0] address_91;
    wire _1505;
    wire read_enable_75;
    wire _1503;
    wire write_enable_91;
    wire _1507;
    wire [131:0] _1515;
    wire [63:0] _1516;
    wire [63:0] _1571;
    wire [63:0] data_87;
    wire [63:0] data_88;
    wire [63:0] data_89;
    wire [63:0] data_90;
    wire [5:0] _198 = 6'b000000;
    wire [5:0] _197 = 6'b000000;
    wire [5:0] _195 = 6'b000000;
    wire [5:0] _194 = 6'b000000;
    wire [5:0] _192 = 6'b000000;
    wire [5:0] _191 = 6'b000000;
    wire [5:0] _189 = 6'b000000;
    wire [5:0] _188 = 6'b000000;
    wire [5:0] _186 = 6'b000000;
    wire [5:0] _185 = 6'b000000;
    wire [5:0] _183 = 6'b000000;
    wire [5:0] _182 = 6'b000000;
    wire [5:0] _180 = 6'b000000;
    wire [5:0] _179 = 6'b000000;
    wire [5:0] _177 = 6'b000000;
    wire [5:0] _176 = 6'b000000;
    wire [5:0] _174 = 6'b000000;
    wire [5:0] _173 = 6'b000000;
    reg [5:0] _175;
    reg [5:0] _178;
    reg [5:0] _181;
    reg [5:0] _184;
    reg [5:0] _187;
    reg [5:0] _190;
    reg [5:0] _193;
    reg [5:0] _196;
    reg [5:0] _199;
    wire [5:0] _172;
    wire [5:0] address_92;
    wire _1496;
    wire read_enable_76;
    wire _1493;
    wire _1494;
    wire write_enable_92;
    wire _1498;
    wire [5:0] address_93;
    wire _1489;
    wire read_enable_77;
    wire _1486;
    wire _1487;
    wire write_enable_93;
    wire _1491;
    wire [131:0] _1501;
    wire [63:0] _1502;
    wire _99;
    wire _1484 = 1'b0;
    wire _1483 = 1'b0;
    wire _1572;
    wire _65;
    reg PHASE_21;
    wire [63:0] q0_6;
    wire _1481 = 1'b0;
    wire _1480 = 1'b0;
    wire _92;
    reg _1482;
    wire [63:0] _1561;
    wire [191:0] _1570;
    wire [63:0] _1573;
    wire [63:0] data_91;
    wire [63:0] data_92;
    wire [63:0] data_93;
    wire [63:0] data_94;
    wire [5:0] _163 = 6'b000000;
    wire [5:0] _162 = 6'b000000;
    wire [5:0] _160 = 6'b000000;
    wire [5:0] _159 = 6'b000000;
    wire [5:0] _157 = 6'b000000;
    wire [5:0] _156 = 6'b000000;
    wire [5:0] _154 = 6'b000000;
    wire [5:0] _153 = 6'b000000;
    wire [5:0] _151 = 6'b000000;
    wire [5:0] _150 = 6'b000000;
    wire [5:0] _148 = 6'b000000;
    wire [5:0] _147 = 6'b000000;
    wire [5:0] _145 = 6'b000000;
    wire [5:0] _144 = 6'b000000;
    wire [5:0] _142 = 6'b000000;
    wire [5:0] _141 = 6'b000000;
    wire [5:0] _139 = 6'b000000;
    wire [5:0] _138 = 6'b000000;
    wire [5:0] _137;
    reg [5:0] _140;
    reg [5:0] _143;
    reg [5:0] _146;
    reg [5:0] _149;
    reg [5:0] _152;
    reg [5:0] _155;
    reg [5:0] _158;
    reg [5:0] _161;
    reg [5:0] _164;
    wire [5:0] _68;
    wire [5:0] address_94;
    wire _1637;
    wire [7:0] _70;
    wire _1636;
    wire read_enable_78;
    wire _1630 = 1'b0;
    wire _1629 = 1'b0;
    wire _1627 = 1'b0;
    wire _1626 = 1'b0;
    wire _1624 = 1'b0;
    wire _1623 = 1'b0;
    wire _1621 = 1'b0;
    wire _1620 = 1'b0;
    wire _1618 = 1'b0;
    wire _1617 = 1'b0;
    wire _1615 = 1'b0;
    wire _1614 = 1'b0;
    wire _1612 = 1'b0;
    wire _1611 = 1'b0;
    wire _1609 = 1'b0;
    wire _1608 = 1'b0;
    wire _1606 = 1'b0;
    wire _1605 = 1'b0;
    wire _278;
    reg _1607;
    reg _1610;
    reg _1613;
    reg _1616;
    reg _1619;
    reg _1622;
    reg _1625;
    reg _1628;
    reg _1631;
    wire _1632;
    wire _1603 = 1'b0;
    wire _1602 = 1'b0;
    wire _1600 = 1'b0;
    wire _1599 = 1'b0;
    wire _1597 = 1'b0;
    wire _1596 = 1'b0;
    wire _1594 = 1'b0;
    wire _1593 = 1'b0;
    wire _1591 = 1'b0;
    wire _1590 = 1'b0;
    wire _1588 = 1'b0;
    wire _1587 = 1'b0;
    wire _1585 = 1'b0;
    wire _1584 = 1'b0;
    wire _1582 = 1'b0;
    wire _1581 = 1'b0;
    wire _1579 = 1'b0;
    wire _1578 = 1'b0;
    wire _130;
    reg _1580;
    reg _1583;
    reg _1586;
    reg _1589;
    reg _1592;
    reg _1595;
    reg _1598;
    reg _1601;
    reg _1604;
    wire _1633;
    wire _128 = 1'b0;
    wire _127 = 1'b0;
    wire _125 = 1'b0;
    wire _124 = 1'b0;
    wire _122 = 1'b0;
    wire _121 = 1'b0;
    wire _119 = 1'b0;
    wire _118 = 1'b0;
    wire _116 = 1'b0;
    wire _115 = 1'b0;
    wire _113 = 1'b0;
    wire _112 = 1'b0;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire vdd = 1'b1;
    wire _104 = 1'b0;
    wire _103 = 1'b0;
    wire _102;
    reg _105;
    reg _108;
    reg _111;
    reg _114;
    reg _117;
    reg _120;
    reg _123;
    reg _126;
    reg _129;
    wire _1634;
    wire write_enable_94;
    wire _1639;
    wire gnd = 1'b0;
    wire [131:0] _1646;
    wire [63:0] _1647;
    wire _72;
    wire _1575 = 1'b0;
    wire _1574 = 1'b0;
    wire _1577;
    wire _73;
    reg PHASE_22;
    wire [63:0] _1659;
    wire _76;
    wire _78;
    wire _80;
    wire _82;
    wire _84;
    wire [492:0] _91;
    wire _1660;

    /* logic */
    assign address = _360 ? _199 : _355;
    assign write_enable = _353 & _360;
    assign address_0 = _360 ? _164 : _68;
    assign _362 = ~ _360;
    assign read_enable = _348 & _362;
    assign _360 = ~ PHASE_1;
    assign write_enable_0 = _346 & _360;
    assign _364 = write_enable_0 | read_enable;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_364), .regcea(vdd), .wea(write_enable_0), .addra(address_0), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable), .regceb(vdd), .web(write_enable), .addrb(address), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_369[131:131]), .sbiterrb(_369[130:130]), .doutb(_369[129:66]), .dbiterra(_369[65:65]), .sbiterra(_369[64:64]), .douta(_369[63:0]) );
    assign _370 = _369[63:0];
    assign address_1 = PHASE_1 ? _199 : _355;
    assign _353 = _129 & _316;
    assign write_enable_1 = _353 & PHASE_1;
    assign _267 = _259[129:66];
    assign _266 = _246[129:66];
    assign _268 = PHASE ? _267 : _266;
    assign _264 = _216[129:66];
    assign _263 = _202[129:66];
    assign q1 = PHASE_0 ? _264 : _263;
    assign _269 = _96 ? _268 : q1;
    assign address_2 = _248 ? _242 : _241;
    assign _254 = ~ _248;
    assign read_enable_0 = _102 & _254;
    assign address_3 = _248 ? _60 : _230;
    assign _250 = ~ _248;
    assign read_enable_1 = _102 & _250;
    assign _248 = ~ PHASE;
    assign write_enable_3 = _219 & _248;
    assign _252 = write_enable_3 | read_enable_1;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_0
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_252), .regcea(vdd), .wea(write_enable_3), .addra(address_3), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_0), .regceb(vdd), .web(write_enable_2), .addrb(address_2), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_259[131:131]), .sbiterrb(_259[130:130]), .doutb(_259[129:66]), .dbiterra(_259[65:65]), .sbiterra(_259[64:64]), .douta(_259[63:0]) );
    assign _260 = _259[63:0];
    assign _240 = _172[5:5];
    assign _239 = _172[4:4];
    assign _238 = _172[3:3];
    assign _237 = _172[2:2];
    assign _236 = _172[1:1];
    assign _235 = _172[0:0];
    assign _241 = { _235, _236, _237, _238, _239, _240 };
    assign address_4 = PHASE ? _242 : _241;
    assign _232 = ~ PHASE;
    assign read_enable_2 = _102 & _232;
    assign data_1 = wr_d7;
    assign _229 = _137[5:5];
    assign _228 = _137[4:4];
    assign _227 = _137[3:3];
    assign _226 = _137[2:2];
    assign _225 = _137[1:1];
    assign _224 = _137[0:0];
    assign _230 = { _224, _225, _226, _227, _228, _229 };
    assign address_5 = PHASE ? _60 : _230;
    assign _221 = ~ PHASE;
    assign read_enable_3 = _102 & _221;
    assign _219 = _62[7:7];
    assign write_enable_5 = _219 & PHASE;
    assign _223 = write_enable_5 | read_enable_3;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_1
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_223), .regcea(vdd), .wea(write_enable_5), .addra(address_5), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_2), .regceb(vdd), .web(write_enable_4), .addrb(address_4), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_246[131:131]), .sbiterrb(_246[130:130]), .doutb(_246[129:66]), .dbiterra(_246[65:65]), .sbiterra(_246[64:64]), .douta(_246[63:0]) );
    assign _247 = _246[63:0];
    assign _89 = ~ PHASE;
    assign _3 = _89;
    always @(posedge _84) begin
        if (_82)
            PHASE <= _87;
        else
            if (_72)
                PHASE <= _3;
    end
    assign _261 = PHASE ? _260 : _247;
    assign address_6 = _204 ? _199 : _172;
    assign _211 = ~ _204;
    assign read_enable_4 = _102 & _211;
    assign write_enable_6 = _167 & _204;
    assign _213 = write_enable_6 | read_enable_4;
    assign address_7 = _204 ? _164 : _137;
    assign _206 = ~ _204;
    assign read_enable_5 = _102 & _206;
    assign _204 = ~ PHASE_0;
    assign write_enable_7 = _132 & _204;
    assign _208 = write_enable_7 | read_enable_5;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_2
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_208), .regcea(vdd), .wea(write_enable_7), .addra(address_7), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_213), .regceb(vdd), .web(write_enable_6), .addrb(address_6), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_216[131:131]), .sbiterrb(_216[130:130]), .doutb(_216[129:66]), .dbiterra(_216[65:65]), .sbiterra(_216[64:64]), .douta(_216[63:0]) );
    assign _217 = _216[63:0];
    assign _283 = _282[127:64];
    assign data_3 = _283;
    assign address_8 = PHASE_0 ? _199 : _172;
    assign _169 = ~ PHASE_0;
    assign read_enable_6 = _102 & _169;
    assign _166 = ~ _130;
    assign _167 = _129 & _166;
    assign write_enable_8 = _167 & PHASE_0;
    assign _171 = write_enable_8 | read_enable_6;
    assign address_9 = PHASE_0 ? _164 : _137;
    assign _134 = ~ PHASE_0;
    assign read_enable_7 = _102 & _134;
    assign _131 = ~ _130;
    assign _132 = _129 & _131;
    assign write_enable_9 = _132 & PHASE_0;
    assign _136 = write_enable_9 | read_enable_7;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_3
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_136), .regcea(vdd), .wea(write_enable_9), .addra(address_9), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_171), .regceb(vdd), .web(write_enable_8), .addrb(address_8), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_202[131:131]), .sbiterrb(_202[130:130]), .doutb(_202[129:66]), .dbiterra(_202[65:65]), .sbiterra(_202[64:64]), .douta(_202[63:0]) );
    assign _203 = _202[63:0];
    assign _284 = ~ PHASE_0;
    assign _5 = _284;
    always @(posedge _84) begin
        if (_82)
            PHASE_0 <= _98;
        else
            if (_99)
                PHASE_0 <= _5;
    end
    assign q0 = PHASE_0 ? _217 : _203;
    always @(posedge _84) begin
        if (_82)
            _96 <= _94;
        else
            _96 <= _92;
    end
    assign _262 = _96 ? _261 : q0;
    dp_6
        dp_6
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_262), .d2(_269), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_282[191:128]), .q2(_282[127:64]), .q1(_282[63:0]) );
    assign _285 = _282[63:0];
    assign data_7 = _285;
    assign address_10 = PHASE_1 ? _164 : _68;
    assign _349 = ~ PHASE_1;
    assign _348 = _70[7:7];
    assign read_enable_8 = _348 & _349;
    always @(posedge _84) begin
        if (_82)
            _319 <= _318;
        else
            _319 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _322 <= _321;
        else
            _322 <= _319;
    end
    always @(posedge _84) begin
        if (_82)
            _325 <= _324;
        else
            _325 <= _322;
    end
    always @(posedge _84) begin
        if (_82)
            _328 <= _327;
        else
            _328 <= _325;
    end
    always @(posedge _84) begin
        if (_82)
            _331 <= _330;
        else
            _331 <= _328;
    end
    always @(posedge _84) begin
        if (_82)
            _334 <= _333;
        else
            _334 <= _331;
    end
    always @(posedge _84) begin
        if (_82)
            _337 <= _336;
        else
            _337 <= _334;
    end
    always @(posedge _84) begin
        if (_82)
            _340 <= _339;
        else
            _340 <= _337;
    end
    always @(posedge _84) begin
        if (_82)
            _343 <= _342;
        else
            _343 <= _340;
    end
    assign _344 = ~ _343;
    always @(posedge _84) begin
        if (_82)
            _292 <= _291;
        else
            _292 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _295 <= _294;
        else
            _295 <= _292;
    end
    always @(posedge _84) begin
        if (_82)
            _298 <= _297;
        else
            _298 <= _295;
    end
    always @(posedge _84) begin
        if (_82)
            _301 <= _300;
        else
            _301 <= _298;
    end
    always @(posedge _84) begin
        if (_82)
            _304 <= _303;
        else
            _304 <= _301;
    end
    always @(posedge _84) begin
        if (_82)
            _307 <= _306;
        else
            _307 <= _304;
    end
    always @(posedge _84) begin
        if (_82)
            _310 <= _309;
        else
            _310 <= _307;
    end
    always @(posedge _84) begin
        if (_82)
            _313 <= _312;
        else
            _313 <= _310;
    end
    always @(posedge _84) begin
        if (_82)
            _316 <= _315;
        else
            _316 <= _313;
    end
    assign _345 = _316 & _344;
    assign _346 = _129 & _345;
    assign write_enable_10 = _346 & PHASE_1;
    assign _351 = write_enable_10 | read_enable_8;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_4
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_351), .regcea(vdd), .wea(write_enable_10), .addra(address_10), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_1), .regceb(vdd), .web(write_enable_1), .addrb(address_1), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_358[131:131]), .sbiterrb(_358[130:130]), .doutb(_358[129:66]), .dbiterra(_358[65:65]), .sbiterra(_358[64:64]), .douta(_358[63:0]) );
    assign _359 = _358[63:0];
    assign _289 = ~ PHASE_1;
    assign _7 = _289;
    always @(posedge _84) begin
        if (_82)
            PHASE_1 <= _287;
        else
            if (_72)
                PHASE_1 <= _7;
    end
    assign _371 = PHASE_1 ? _370 : _359;
    assign address_11 = _544 ? _199 : _539;
    assign write_enable_11 = _537 & _544;
    assign address_12 = _544 ? _164 : _68;
    assign _546 = ~ _544;
    assign read_enable_9 = _532 & _546;
    assign _544 = ~ PHASE_4;
    assign write_enable_12 = _530 & _544;
    assign _548 = write_enable_12 | read_enable_9;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_5
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_548), .regcea(vdd), .wea(write_enable_12), .addra(address_12), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_11), .regceb(vdd), .web(write_enable_11), .addrb(address_11), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_553[131:131]), .sbiterrb(_553[130:130]), .doutb(_553[129:66]), .dbiterra(_553[65:65]), .sbiterra(_553[64:64]), .douta(_553[63:0]) );
    assign _554 = _553[63:0];
    assign address_13 = PHASE_4 ? _199 : _539;
    assign _537 = _129 & _500;
    assign write_enable_13 = _537 & PHASE_4;
    assign _462 = _454[129:66];
    assign _461 = _441[129:66];
    assign _463 = PHASE_2 ? _462 : _461;
    assign _459 = _411[129:66];
    assign _458 = _397[129:66];
    assign q1_0 = PHASE_3 ? _459 : _458;
    assign _464 = _378 ? _463 : q1_0;
    assign address_14 = _443 ? _437 : _436;
    assign _449 = ~ _443;
    assign read_enable_10 = _102 & _449;
    assign address_15 = _443 ? _60 : _425;
    assign _445 = ~ _443;
    assign read_enable_11 = _102 & _445;
    assign _443 = ~ PHASE_2;
    assign write_enable_15 = _414 & _443;
    assign _447 = write_enable_15 | read_enable_11;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_6
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_447), .regcea(vdd), .wea(write_enable_15), .addra(address_15), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_10), .regceb(vdd), .web(write_enable_14), .addrb(address_14), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_454[131:131]), .sbiterrb(_454[130:130]), .doutb(_454[129:66]), .dbiterra(_454[65:65]), .sbiterra(_454[64:64]), .douta(_454[63:0]) );
    assign _455 = _454[63:0];
    assign _435 = _172[5:5];
    assign _434 = _172[4:4];
    assign _433 = _172[3:3];
    assign _432 = _172[2:2];
    assign _431 = _172[1:1];
    assign _430 = _172[0:0];
    assign _436 = { _430, _431, _432, _433, _434, _435 };
    assign address_16 = PHASE_2 ? _437 : _436;
    assign _427 = ~ PHASE_2;
    assign read_enable_12 = _102 & _427;
    assign data_13 = wr_d6;
    assign _424 = _137[5:5];
    assign _423 = _137[4:4];
    assign _422 = _137[3:3];
    assign _421 = _137[2:2];
    assign _420 = _137[1:1];
    assign _419 = _137[0:0];
    assign _425 = { _419, _420, _421, _422, _423, _424 };
    assign address_17 = PHASE_2 ? _60 : _425;
    assign _416 = ~ PHASE_2;
    assign read_enable_13 = _102 & _416;
    assign _414 = _62[6:6];
    assign write_enable_17 = _414 & PHASE_2;
    assign _418 = write_enable_17 | read_enable_13;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_7
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_418), .regcea(vdd), .wea(write_enable_17), .addra(address_17), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_12), .regceb(vdd), .web(write_enable_16), .addrb(address_16), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_441[131:131]), .sbiterrb(_441[130:130]), .doutb(_441[129:66]), .dbiterra(_441[65:65]), .sbiterra(_441[64:64]), .douta(_441[63:0]) );
    assign _442 = _441[63:0];
    assign _375 = ~ PHASE_2;
    assign _11 = _375;
    always @(posedge _84) begin
        if (_82)
            PHASE_2 <= _373;
        else
            if (_72)
                PHASE_2 <= _11;
    end
    assign _456 = PHASE_2 ? _455 : _442;
    assign address_18 = _399 ? _199 : _172;
    assign _406 = ~ _399;
    assign read_enable_14 = _102 & _406;
    assign write_enable_18 = _390 & _399;
    assign _408 = write_enable_18 | read_enable_14;
    assign address_19 = _399 ? _164 : _137;
    assign _401 = ~ _399;
    assign read_enable_15 = _102 & _401;
    assign _399 = ~ PHASE_3;
    assign write_enable_19 = _383 & _399;
    assign _403 = write_enable_19 | read_enable_15;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_8
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_403), .regcea(vdd), .wea(write_enable_19), .addra(address_19), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_408), .regceb(vdd), .web(write_enable_18), .addrb(address_18), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_411[131:131]), .sbiterrb(_411[130:130]), .doutb(_411[129:66]), .dbiterra(_411[65:65]), .sbiterra(_411[64:64]), .douta(_411[63:0]) );
    assign _412 = _411[63:0];
    assign _467 = _466[127:64];
    assign data_15 = _467;
    assign address_20 = PHASE_3 ? _199 : _172;
    assign _392 = ~ PHASE_3;
    assign read_enable_16 = _102 & _392;
    assign _389 = ~ _130;
    assign _390 = _129 & _389;
    assign write_enable_20 = _390 & PHASE_3;
    assign _394 = write_enable_20 | read_enable_16;
    assign address_21 = PHASE_3 ? _164 : _137;
    assign _385 = ~ PHASE_3;
    assign read_enable_17 = _102 & _385;
    assign _382 = ~ _130;
    assign _383 = _129 & _382;
    assign write_enable_21 = _383 & PHASE_3;
    assign _387 = write_enable_21 | read_enable_17;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_9
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_387), .regcea(vdd), .wea(write_enable_21), .addra(address_21), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_394), .regceb(vdd), .web(write_enable_20), .addrb(address_20), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_397[131:131]), .sbiterrb(_397[130:130]), .doutb(_397[129:66]), .dbiterra(_397[65:65]), .sbiterra(_397[64:64]), .douta(_397[63:0]) );
    assign _398 = _397[63:0];
    assign _468 = ~ PHASE_3;
    assign _13 = _468;
    always @(posedge _84) begin
        if (_82)
            PHASE_3 <= _380;
        else
            if (_99)
                PHASE_3 <= _13;
    end
    assign q0_0 = PHASE_3 ? _412 : _398;
    always @(posedge _84) begin
        if (_82)
            _378 <= _377;
        else
            _378 <= _92;
    end
    assign _457 = _378 ? _456 : q0_0;
    dp_5
        dp_5
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_457), .d2(_464), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_466[191:128]), .q2(_466[127:64]), .q1(_466[63:0]) );
    assign _469 = _466[63:0];
    assign data_19 = _469;
    assign address_22 = PHASE_4 ? _164 : _68;
    assign _533 = ~ PHASE_4;
    assign _532 = _70[6:6];
    assign read_enable_18 = _532 & _533;
    always @(posedge _84) begin
        if (_82)
            _503 <= _502;
        else
            _503 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _506 <= _505;
        else
            _506 <= _503;
    end
    always @(posedge _84) begin
        if (_82)
            _509 <= _508;
        else
            _509 <= _506;
    end
    always @(posedge _84) begin
        if (_82)
            _512 <= _511;
        else
            _512 <= _509;
    end
    always @(posedge _84) begin
        if (_82)
            _515 <= _514;
        else
            _515 <= _512;
    end
    always @(posedge _84) begin
        if (_82)
            _518 <= _517;
        else
            _518 <= _515;
    end
    always @(posedge _84) begin
        if (_82)
            _521 <= _520;
        else
            _521 <= _518;
    end
    always @(posedge _84) begin
        if (_82)
            _524 <= _523;
        else
            _524 <= _521;
    end
    always @(posedge _84) begin
        if (_82)
            _527 <= _526;
        else
            _527 <= _524;
    end
    assign _528 = ~ _527;
    always @(posedge _84) begin
        if (_82)
            _476 <= _475;
        else
            _476 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _479 <= _478;
        else
            _479 <= _476;
    end
    always @(posedge _84) begin
        if (_82)
            _482 <= _481;
        else
            _482 <= _479;
    end
    always @(posedge _84) begin
        if (_82)
            _485 <= _484;
        else
            _485 <= _482;
    end
    always @(posedge _84) begin
        if (_82)
            _488 <= _487;
        else
            _488 <= _485;
    end
    always @(posedge _84) begin
        if (_82)
            _491 <= _490;
        else
            _491 <= _488;
    end
    always @(posedge _84) begin
        if (_82)
            _494 <= _493;
        else
            _494 <= _491;
    end
    always @(posedge _84) begin
        if (_82)
            _497 <= _496;
        else
            _497 <= _494;
    end
    always @(posedge _84) begin
        if (_82)
            _500 <= _499;
        else
            _500 <= _497;
    end
    assign _529 = _500 & _528;
    assign _530 = _129 & _529;
    assign write_enable_22 = _530 & PHASE_4;
    assign _535 = write_enable_22 | read_enable_18;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_10
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_535), .regcea(vdd), .wea(write_enable_22), .addra(address_22), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_13), .regceb(vdd), .web(write_enable_13), .addrb(address_13), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_542[131:131]), .sbiterrb(_542[130:130]), .doutb(_542[129:66]), .dbiterra(_542[65:65]), .sbiterra(_542[64:64]), .douta(_542[63:0]) );
    assign _543 = _542[63:0];
    assign _473 = ~ PHASE_4;
    assign _15 = _473;
    always @(posedge _84) begin
        if (_82)
            PHASE_4 <= _471;
        else
            if (_72)
                PHASE_4 <= _15;
    end
    assign _555 = PHASE_4 ? _554 : _543;
    assign address_23 = _728 ? _199 : _723;
    assign write_enable_23 = _721 & _728;
    assign address_24 = _728 ? _164 : _68;
    assign _730 = ~ _728;
    assign read_enable_19 = _716 & _730;
    assign _728 = ~ PHASE_7;
    assign write_enable_24 = _714 & _728;
    assign _732 = write_enable_24 | read_enable_19;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_11
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_732), .regcea(vdd), .wea(write_enable_24), .addra(address_24), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_23), .regceb(vdd), .web(write_enable_23), .addrb(address_23), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_737[131:131]), .sbiterrb(_737[130:130]), .doutb(_737[129:66]), .dbiterra(_737[65:65]), .sbiterra(_737[64:64]), .douta(_737[63:0]) );
    assign _738 = _737[63:0];
    assign address_25 = PHASE_7 ? _199 : _723;
    assign _721 = _129 & _684;
    assign write_enable_25 = _721 & PHASE_7;
    assign _646 = _638[129:66];
    assign _645 = _625[129:66];
    assign _647 = PHASE_5 ? _646 : _645;
    assign _643 = _595[129:66];
    assign _642 = _581[129:66];
    assign q1_1 = PHASE_6 ? _643 : _642;
    assign _648 = _562 ? _647 : q1_1;
    assign address_26 = _627 ? _621 : _620;
    assign _633 = ~ _627;
    assign read_enable_20 = _102 & _633;
    assign address_27 = _627 ? _60 : _609;
    assign _629 = ~ _627;
    assign read_enable_21 = _102 & _629;
    assign _627 = ~ PHASE_5;
    assign write_enable_27 = _598 & _627;
    assign _631 = write_enable_27 | read_enable_21;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_12
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_631), .regcea(vdd), .wea(write_enable_27), .addra(address_27), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_20), .regceb(vdd), .web(write_enable_26), .addrb(address_26), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_638[131:131]), .sbiterrb(_638[130:130]), .doutb(_638[129:66]), .dbiterra(_638[65:65]), .sbiterra(_638[64:64]), .douta(_638[63:0]) );
    assign _639 = _638[63:0];
    assign _619 = _172[5:5];
    assign _618 = _172[4:4];
    assign _617 = _172[3:3];
    assign _616 = _172[2:2];
    assign _615 = _172[1:1];
    assign _614 = _172[0:0];
    assign _620 = { _614, _615, _616, _617, _618, _619 };
    assign address_28 = PHASE_5 ? _621 : _620;
    assign _611 = ~ PHASE_5;
    assign read_enable_22 = _102 & _611;
    assign data_25 = wr_d5;
    assign _608 = _137[5:5];
    assign _607 = _137[4:4];
    assign _606 = _137[3:3];
    assign _605 = _137[2:2];
    assign _604 = _137[1:1];
    assign _603 = _137[0:0];
    assign _609 = { _603, _604, _605, _606, _607, _608 };
    assign address_29 = PHASE_5 ? _60 : _609;
    assign _600 = ~ PHASE_5;
    assign read_enable_23 = _102 & _600;
    assign _598 = _62[5:5];
    assign write_enable_29 = _598 & PHASE_5;
    assign _602 = write_enable_29 | read_enable_23;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_13
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_602), .regcea(vdd), .wea(write_enable_29), .addra(address_29), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_22), .regceb(vdd), .web(write_enable_28), .addrb(address_28), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_625[131:131]), .sbiterrb(_625[130:130]), .doutb(_625[129:66]), .dbiterra(_625[65:65]), .sbiterra(_625[64:64]), .douta(_625[63:0]) );
    assign _626 = _625[63:0];
    assign _559 = ~ PHASE_5;
    assign _19 = _559;
    always @(posedge _84) begin
        if (_82)
            PHASE_5 <= _557;
        else
            if (_72)
                PHASE_5 <= _19;
    end
    assign _640 = PHASE_5 ? _639 : _626;
    assign address_30 = _583 ? _199 : _172;
    assign _590 = ~ _583;
    assign read_enable_24 = _102 & _590;
    assign write_enable_30 = _574 & _583;
    assign _592 = write_enable_30 | read_enable_24;
    assign address_31 = _583 ? _164 : _137;
    assign _585 = ~ _583;
    assign read_enable_25 = _102 & _585;
    assign _583 = ~ PHASE_6;
    assign write_enable_31 = _567 & _583;
    assign _587 = write_enable_31 | read_enable_25;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_14
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_587), .regcea(vdd), .wea(write_enable_31), .addra(address_31), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_592), .regceb(vdd), .web(write_enable_30), .addrb(address_30), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_595[131:131]), .sbiterrb(_595[130:130]), .doutb(_595[129:66]), .dbiterra(_595[65:65]), .sbiterra(_595[64:64]), .douta(_595[63:0]) );
    assign _596 = _595[63:0];
    assign _651 = _650[127:64];
    assign data_27 = _651;
    assign address_32 = PHASE_6 ? _199 : _172;
    assign _576 = ~ PHASE_6;
    assign read_enable_26 = _102 & _576;
    assign _573 = ~ _130;
    assign _574 = _129 & _573;
    assign write_enable_32 = _574 & PHASE_6;
    assign _578 = write_enable_32 | read_enable_26;
    assign address_33 = PHASE_6 ? _164 : _137;
    assign _569 = ~ PHASE_6;
    assign read_enable_27 = _102 & _569;
    assign _566 = ~ _130;
    assign _567 = _129 & _566;
    assign write_enable_33 = _567 & PHASE_6;
    assign _571 = write_enable_33 | read_enable_27;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_15
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_571), .regcea(vdd), .wea(write_enable_33), .addra(address_33), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_578), .regceb(vdd), .web(write_enable_32), .addrb(address_32), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_581[131:131]), .sbiterrb(_581[130:130]), .doutb(_581[129:66]), .dbiterra(_581[65:65]), .sbiterra(_581[64:64]), .douta(_581[63:0]) );
    assign _582 = _581[63:0];
    assign _652 = ~ PHASE_6;
    assign _21 = _652;
    always @(posedge _84) begin
        if (_82)
            PHASE_6 <= _564;
        else
            if (_99)
                PHASE_6 <= _21;
    end
    assign q0_1 = PHASE_6 ? _596 : _582;
    always @(posedge _84) begin
        if (_82)
            _562 <= _561;
        else
            _562 <= _92;
    end
    assign _641 = _562 ? _640 : q0_1;
    dp_4
        dp_4
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_641), .d2(_648), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_650[191:128]), .q2(_650[127:64]), .q1(_650[63:0]) );
    assign _653 = _650[63:0];
    assign data_31 = _653;
    assign address_34 = PHASE_7 ? _164 : _68;
    assign _717 = ~ PHASE_7;
    assign _716 = _70[5:5];
    assign read_enable_28 = _716 & _717;
    always @(posedge _84) begin
        if (_82)
            _687 <= _686;
        else
            _687 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _690 <= _689;
        else
            _690 <= _687;
    end
    always @(posedge _84) begin
        if (_82)
            _693 <= _692;
        else
            _693 <= _690;
    end
    always @(posedge _84) begin
        if (_82)
            _696 <= _695;
        else
            _696 <= _693;
    end
    always @(posedge _84) begin
        if (_82)
            _699 <= _698;
        else
            _699 <= _696;
    end
    always @(posedge _84) begin
        if (_82)
            _702 <= _701;
        else
            _702 <= _699;
    end
    always @(posedge _84) begin
        if (_82)
            _705 <= _704;
        else
            _705 <= _702;
    end
    always @(posedge _84) begin
        if (_82)
            _708 <= _707;
        else
            _708 <= _705;
    end
    always @(posedge _84) begin
        if (_82)
            _711 <= _710;
        else
            _711 <= _708;
    end
    assign _712 = ~ _711;
    always @(posedge _84) begin
        if (_82)
            _660 <= _659;
        else
            _660 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _663 <= _662;
        else
            _663 <= _660;
    end
    always @(posedge _84) begin
        if (_82)
            _666 <= _665;
        else
            _666 <= _663;
    end
    always @(posedge _84) begin
        if (_82)
            _669 <= _668;
        else
            _669 <= _666;
    end
    always @(posedge _84) begin
        if (_82)
            _672 <= _671;
        else
            _672 <= _669;
    end
    always @(posedge _84) begin
        if (_82)
            _675 <= _674;
        else
            _675 <= _672;
    end
    always @(posedge _84) begin
        if (_82)
            _678 <= _677;
        else
            _678 <= _675;
    end
    always @(posedge _84) begin
        if (_82)
            _681 <= _680;
        else
            _681 <= _678;
    end
    always @(posedge _84) begin
        if (_82)
            _684 <= _683;
        else
            _684 <= _681;
    end
    assign _713 = _684 & _712;
    assign _714 = _129 & _713;
    assign write_enable_34 = _714 & PHASE_7;
    assign _719 = write_enable_34 | read_enable_28;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_16
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_719), .regcea(vdd), .wea(write_enable_34), .addra(address_34), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_25), .regceb(vdd), .web(write_enable_25), .addrb(address_25), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_726[131:131]), .sbiterrb(_726[130:130]), .doutb(_726[129:66]), .dbiterra(_726[65:65]), .sbiterra(_726[64:64]), .douta(_726[63:0]) );
    assign _727 = _726[63:0];
    assign _657 = ~ PHASE_7;
    assign _23 = _657;
    always @(posedge _84) begin
        if (_82)
            PHASE_7 <= _655;
        else
            if (_72)
                PHASE_7 <= _23;
    end
    assign _739 = PHASE_7 ? _738 : _727;
    assign address_35 = _912 ? _199 : _907;
    assign write_enable_35 = _905 & _912;
    assign address_36 = _912 ? _164 : _68;
    assign _914 = ~ _912;
    assign read_enable_29 = _900 & _914;
    assign _912 = ~ PHASE_10;
    assign write_enable_36 = _898 & _912;
    assign _916 = write_enable_36 | read_enable_29;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_17
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_916), .regcea(vdd), .wea(write_enable_36), .addra(address_36), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_35), .regceb(vdd), .web(write_enable_35), .addrb(address_35), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_921[131:131]), .sbiterrb(_921[130:130]), .doutb(_921[129:66]), .dbiterra(_921[65:65]), .sbiterra(_921[64:64]), .douta(_921[63:0]) );
    assign _922 = _921[63:0];
    assign address_37 = PHASE_10 ? _199 : _907;
    assign _905 = _129 & _868;
    assign write_enable_37 = _905 & PHASE_10;
    assign _830 = _822[129:66];
    assign _829 = _809[129:66];
    assign _831 = PHASE_8 ? _830 : _829;
    assign _827 = _779[129:66];
    assign _826 = _765[129:66];
    assign q1_2 = PHASE_9 ? _827 : _826;
    assign _832 = _746 ? _831 : q1_2;
    assign address_38 = _811 ? _805 : _804;
    assign _817 = ~ _811;
    assign read_enable_30 = _102 & _817;
    assign address_39 = _811 ? _60 : _793;
    assign _813 = ~ _811;
    assign read_enable_31 = _102 & _813;
    assign _811 = ~ PHASE_8;
    assign write_enable_39 = _782 & _811;
    assign _815 = write_enable_39 | read_enable_31;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_18
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_815), .regcea(vdd), .wea(write_enable_39), .addra(address_39), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_30), .regceb(vdd), .web(write_enable_38), .addrb(address_38), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_822[131:131]), .sbiterrb(_822[130:130]), .doutb(_822[129:66]), .dbiterra(_822[65:65]), .sbiterra(_822[64:64]), .douta(_822[63:0]) );
    assign _823 = _822[63:0];
    assign _803 = _172[5:5];
    assign _802 = _172[4:4];
    assign _801 = _172[3:3];
    assign _800 = _172[2:2];
    assign _799 = _172[1:1];
    assign _798 = _172[0:0];
    assign _804 = { _798, _799, _800, _801, _802, _803 };
    assign address_40 = PHASE_8 ? _805 : _804;
    assign _795 = ~ PHASE_8;
    assign read_enable_32 = _102 & _795;
    assign data_37 = wr_d4;
    assign _792 = _137[5:5];
    assign _791 = _137[4:4];
    assign _790 = _137[3:3];
    assign _789 = _137[2:2];
    assign _788 = _137[1:1];
    assign _787 = _137[0:0];
    assign _793 = { _787, _788, _789, _790, _791, _792 };
    assign address_41 = PHASE_8 ? _60 : _793;
    assign _784 = ~ PHASE_8;
    assign read_enable_33 = _102 & _784;
    assign _782 = _62[4:4];
    assign write_enable_41 = _782 & PHASE_8;
    assign _786 = write_enable_41 | read_enable_33;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_19
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_786), .regcea(vdd), .wea(write_enable_41), .addra(address_41), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_32), .regceb(vdd), .web(write_enable_40), .addrb(address_40), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_809[131:131]), .sbiterrb(_809[130:130]), .doutb(_809[129:66]), .dbiterra(_809[65:65]), .sbiterra(_809[64:64]), .douta(_809[63:0]) );
    assign _810 = _809[63:0];
    assign _743 = ~ PHASE_8;
    assign _27 = _743;
    always @(posedge _84) begin
        if (_82)
            PHASE_8 <= _741;
        else
            if (_72)
                PHASE_8 <= _27;
    end
    assign _824 = PHASE_8 ? _823 : _810;
    assign address_42 = _767 ? _199 : _172;
    assign _774 = ~ _767;
    assign read_enable_34 = _102 & _774;
    assign write_enable_42 = _758 & _767;
    assign _776 = write_enable_42 | read_enable_34;
    assign address_43 = _767 ? _164 : _137;
    assign _769 = ~ _767;
    assign read_enable_35 = _102 & _769;
    assign _767 = ~ PHASE_9;
    assign write_enable_43 = _751 & _767;
    assign _771 = write_enable_43 | read_enable_35;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_20
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_771), .regcea(vdd), .wea(write_enable_43), .addra(address_43), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_776), .regceb(vdd), .web(write_enable_42), .addrb(address_42), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_779[131:131]), .sbiterrb(_779[130:130]), .doutb(_779[129:66]), .dbiterra(_779[65:65]), .sbiterra(_779[64:64]), .douta(_779[63:0]) );
    assign _780 = _779[63:0];
    assign _835 = _834[127:64];
    assign data_39 = _835;
    assign address_44 = PHASE_9 ? _199 : _172;
    assign _760 = ~ PHASE_9;
    assign read_enable_36 = _102 & _760;
    assign _757 = ~ _130;
    assign _758 = _129 & _757;
    assign write_enable_44 = _758 & PHASE_9;
    assign _762 = write_enable_44 | read_enable_36;
    assign address_45 = PHASE_9 ? _164 : _137;
    assign _753 = ~ PHASE_9;
    assign read_enable_37 = _102 & _753;
    assign _750 = ~ _130;
    assign _751 = _129 & _750;
    assign write_enable_45 = _751 & PHASE_9;
    assign _755 = write_enable_45 | read_enable_37;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_21
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_755), .regcea(vdd), .wea(write_enable_45), .addra(address_45), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_762), .regceb(vdd), .web(write_enable_44), .addrb(address_44), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_765[131:131]), .sbiterrb(_765[130:130]), .doutb(_765[129:66]), .dbiterra(_765[65:65]), .sbiterra(_765[64:64]), .douta(_765[63:0]) );
    assign _766 = _765[63:0];
    assign _836 = ~ PHASE_9;
    assign _29 = _836;
    always @(posedge _84) begin
        if (_82)
            PHASE_9 <= _748;
        else
            if (_99)
                PHASE_9 <= _29;
    end
    assign q0_2 = PHASE_9 ? _780 : _766;
    always @(posedge _84) begin
        if (_82)
            _746 <= _745;
        else
            _746 <= _92;
    end
    assign _825 = _746 ? _824 : q0_2;
    dp_3
        dp_3
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_825), .d2(_832), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_834[191:128]), .q2(_834[127:64]), .q1(_834[63:0]) );
    assign _837 = _834[63:0];
    assign data_43 = _837;
    assign address_46 = PHASE_10 ? _164 : _68;
    assign _901 = ~ PHASE_10;
    assign _900 = _70[4:4];
    assign read_enable_38 = _900 & _901;
    always @(posedge _84) begin
        if (_82)
            _871 <= _870;
        else
            _871 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _874 <= _873;
        else
            _874 <= _871;
    end
    always @(posedge _84) begin
        if (_82)
            _877 <= _876;
        else
            _877 <= _874;
    end
    always @(posedge _84) begin
        if (_82)
            _880 <= _879;
        else
            _880 <= _877;
    end
    always @(posedge _84) begin
        if (_82)
            _883 <= _882;
        else
            _883 <= _880;
    end
    always @(posedge _84) begin
        if (_82)
            _886 <= _885;
        else
            _886 <= _883;
    end
    always @(posedge _84) begin
        if (_82)
            _889 <= _888;
        else
            _889 <= _886;
    end
    always @(posedge _84) begin
        if (_82)
            _892 <= _891;
        else
            _892 <= _889;
    end
    always @(posedge _84) begin
        if (_82)
            _895 <= _894;
        else
            _895 <= _892;
    end
    assign _896 = ~ _895;
    always @(posedge _84) begin
        if (_82)
            _844 <= _843;
        else
            _844 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _847 <= _846;
        else
            _847 <= _844;
    end
    always @(posedge _84) begin
        if (_82)
            _850 <= _849;
        else
            _850 <= _847;
    end
    always @(posedge _84) begin
        if (_82)
            _853 <= _852;
        else
            _853 <= _850;
    end
    always @(posedge _84) begin
        if (_82)
            _856 <= _855;
        else
            _856 <= _853;
    end
    always @(posedge _84) begin
        if (_82)
            _859 <= _858;
        else
            _859 <= _856;
    end
    always @(posedge _84) begin
        if (_82)
            _862 <= _861;
        else
            _862 <= _859;
    end
    always @(posedge _84) begin
        if (_82)
            _865 <= _864;
        else
            _865 <= _862;
    end
    always @(posedge _84) begin
        if (_82)
            _868 <= _867;
        else
            _868 <= _865;
    end
    assign _897 = _868 & _896;
    assign _898 = _129 & _897;
    assign write_enable_46 = _898 & PHASE_10;
    assign _903 = write_enable_46 | read_enable_38;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_22
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_903), .regcea(vdd), .wea(write_enable_46), .addra(address_46), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_37), .regceb(vdd), .web(write_enable_37), .addrb(address_37), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_910[131:131]), .sbiterrb(_910[130:130]), .doutb(_910[129:66]), .dbiterra(_910[65:65]), .sbiterra(_910[64:64]), .douta(_910[63:0]) );
    assign _911 = _910[63:0];
    assign _841 = ~ PHASE_10;
    assign _31 = _841;
    always @(posedge _84) begin
        if (_82)
            PHASE_10 <= _839;
        else
            if (_72)
                PHASE_10 <= _31;
    end
    assign _923 = PHASE_10 ? _922 : _911;
    assign address_47 = _1096 ? _199 : _1091;
    assign write_enable_47 = _1089 & _1096;
    assign address_48 = _1096 ? _164 : _68;
    assign _1098 = ~ _1096;
    assign read_enable_39 = _1084 & _1098;
    assign _1096 = ~ PHASE_13;
    assign write_enable_48 = _1082 & _1096;
    assign _1100 = write_enable_48 | read_enable_39;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_23
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1100), .regcea(vdd), .wea(write_enable_48), .addra(address_48), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_47), .regceb(vdd), .web(write_enable_47), .addrb(address_47), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1105[131:131]), .sbiterrb(_1105[130:130]), .doutb(_1105[129:66]), .dbiterra(_1105[65:65]), .sbiterra(_1105[64:64]), .douta(_1105[63:0]) );
    assign _1106 = _1105[63:0];
    assign address_49 = PHASE_13 ? _199 : _1091;
    assign _1089 = _129 & _1052;
    assign write_enable_49 = _1089 & PHASE_13;
    assign _1014 = _1006[129:66];
    assign _1013 = _993[129:66];
    assign _1015 = PHASE_11 ? _1014 : _1013;
    assign _1011 = _963[129:66];
    assign _1010 = _949[129:66];
    assign q1_3 = PHASE_12 ? _1011 : _1010;
    assign _1016 = _930 ? _1015 : q1_3;
    assign address_50 = _995 ? _989 : _988;
    assign _1001 = ~ _995;
    assign read_enable_40 = _102 & _1001;
    assign address_51 = _995 ? _60 : _977;
    assign _997 = ~ _995;
    assign read_enable_41 = _102 & _997;
    assign _995 = ~ PHASE_11;
    assign write_enable_51 = _966 & _995;
    assign _999 = write_enable_51 | read_enable_41;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_24
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_999), .regcea(vdd), .wea(write_enable_51), .addra(address_51), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_40), .regceb(vdd), .web(write_enable_50), .addrb(address_50), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1006[131:131]), .sbiterrb(_1006[130:130]), .doutb(_1006[129:66]), .dbiterra(_1006[65:65]), .sbiterra(_1006[64:64]), .douta(_1006[63:0]) );
    assign _1007 = _1006[63:0];
    assign _987 = _172[5:5];
    assign _986 = _172[4:4];
    assign _985 = _172[3:3];
    assign _984 = _172[2:2];
    assign _983 = _172[1:1];
    assign _982 = _172[0:0];
    assign _988 = { _982, _983, _984, _985, _986, _987 };
    assign address_52 = PHASE_11 ? _989 : _988;
    assign _979 = ~ PHASE_11;
    assign read_enable_42 = _102 & _979;
    assign data_49 = wr_d3;
    assign _976 = _137[5:5];
    assign _975 = _137[4:4];
    assign _974 = _137[3:3];
    assign _973 = _137[2:2];
    assign _972 = _137[1:1];
    assign _971 = _137[0:0];
    assign _977 = { _971, _972, _973, _974, _975, _976 };
    assign address_53 = PHASE_11 ? _60 : _977;
    assign _968 = ~ PHASE_11;
    assign read_enable_43 = _102 & _968;
    assign _966 = _62[3:3];
    assign write_enable_53 = _966 & PHASE_11;
    assign _970 = write_enable_53 | read_enable_43;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_25
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_970), .regcea(vdd), .wea(write_enable_53), .addra(address_53), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_42), .regceb(vdd), .web(write_enable_52), .addrb(address_52), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_993[131:131]), .sbiterrb(_993[130:130]), .doutb(_993[129:66]), .dbiterra(_993[65:65]), .sbiterra(_993[64:64]), .douta(_993[63:0]) );
    assign _994 = _993[63:0];
    assign _927 = ~ PHASE_11;
    assign _35 = _927;
    always @(posedge _84) begin
        if (_82)
            PHASE_11 <= _925;
        else
            if (_72)
                PHASE_11 <= _35;
    end
    assign _1008 = PHASE_11 ? _1007 : _994;
    assign address_54 = _951 ? _199 : _172;
    assign _958 = ~ _951;
    assign read_enable_44 = _102 & _958;
    assign write_enable_54 = _942 & _951;
    assign _960 = write_enable_54 | read_enable_44;
    assign address_55 = _951 ? _164 : _137;
    assign _953 = ~ _951;
    assign read_enable_45 = _102 & _953;
    assign _951 = ~ PHASE_12;
    assign write_enable_55 = _935 & _951;
    assign _955 = write_enable_55 | read_enable_45;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_26
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_955), .regcea(vdd), .wea(write_enable_55), .addra(address_55), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_960), .regceb(vdd), .web(write_enable_54), .addrb(address_54), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_963[131:131]), .sbiterrb(_963[130:130]), .doutb(_963[129:66]), .dbiterra(_963[65:65]), .sbiterra(_963[64:64]), .douta(_963[63:0]) );
    assign _964 = _963[63:0];
    assign _1019 = _1018[127:64];
    assign data_51 = _1019;
    assign address_56 = PHASE_12 ? _199 : _172;
    assign _944 = ~ PHASE_12;
    assign read_enable_46 = _102 & _944;
    assign _941 = ~ _130;
    assign _942 = _129 & _941;
    assign write_enable_56 = _942 & PHASE_12;
    assign _946 = write_enable_56 | read_enable_46;
    assign address_57 = PHASE_12 ? _164 : _137;
    assign _937 = ~ PHASE_12;
    assign read_enable_47 = _102 & _937;
    assign _934 = ~ _130;
    assign _935 = _129 & _934;
    assign write_enable_57 = _935 & PHASE_12;
    assign _939 = write_enable_57 | read_enable_47;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_27
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_939), .regcea(vdd), .wea(write_enable_57), .addra(address_57), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_946), .regceb(vdd), .web(write_enable_56), .addrb(address_56), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_949[131:131]), .sbiterrb(_949[130:130]), .doutb(_949[129:66]), .dbiterra(_949[65:65]), .sbiterra(_949[64:64]), .douta(_949[63:0]) );
    assign _950 = _949[63:0];
    assign _1020 = ~ PHASE_12;
    assign _37 = _1020;
    always @(posedge _84) begin
        if (_82)
            PHASE_12 <= _932;
        else
            if (_99)
                PHASE_12 <= _37;
    end
    assign q0_3 = PHASE_12 ? _964 : _950;
    always @(posedge _84) begin
        if (_82)
            _930 <= _929;
        else
            _930 <= _92;
    end
    assign _1009 = _930 ? _1008 : q0_3;
    dp_2
        dp_2
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1009), .d2(_1016), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_1018[191:128]), .q2(_1018[127:64]), .q1(_1018[63:0]) );
    assign _1021 = _1018[63:0];
    assign data_55 = _1021;
    assign address_58 = PHASE_13 ? _164 : _68;
    assign _1085 = ~ PHASE_13;
    assign _1084 = _70[3:3];
    assign read_enable_48 = _1084 & _1085;
    always @(posedge _84) begin
        if (_82)
            _1055 <= _1054;
        else
            _1055 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _1058 <= _1057;
        else
            _1058 <= _1055;
    end
    always @(posedge _84) begin
        if (_82)
            _1061 <= _1060;
        else
            _1061 <= _1058;
    end
    always @(posedge _84) begin
        if (_82)
            _1064 <= _1063;
        else
            _1064 <= _1061;
    end
    always @(posedge _84) begin
        if (_82)
            _1067 <= _1066;
        else
            _1067 <= _1064;
    end
    always @(posedge _84) begin
        if (_82)
            _1070 <= _1069;
        else
            _1070 <= _1067;
    end
    always @(posedge _84) begin
        if (_82)
            _1073 <= _1072;
        else
            _1073 <= _1070;
    end
    always @(posedge _84) begin
        if (_82)
            _1076 <= _1075;
        else
            _1076 <= _1073;
    end
    always @(posedge _84) begin
        if (_82)
            _1079 <= _1078;
        else
            _1079 <= _1076;
    end
    assign _1080 = ~ _1079;
    always @(posedge _84) begin
        if (_82)
            _1028 <= _1027;
        else
            _1028 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1031 <= _1030;
        else
            _1031 <= _1028;
    end
    always @(posedge _84) begin
        if (_82)
            _1034 <= _1033;
        else
            _1034 <= _1031;
    end
    always @(posedge _84) begin
        if (_82)
            _1037 <= _1036;
        else
            _1037 <= _1034;
    end
    always @(posedge _84) begin
        if (_82)
            _1040 <= _1039;
        else
            _1040 <= _1037;
    end
    always @(posedge _84) begin
        if (_82)
            _1043 <= _1042;
        else
            _1043 <= _1040;
    end
    always @(posedge _84) begin
        if (_82)
            _1046 <= _1045;
        else
            _1046 <= _1043;
    end
    always @(posedge _84) begin
        if (_82)
            _1049 <= _1048;
        else
            _1049 <= _1046;
    end
    always @(posedge _84) begin
        if (_82)
            _1052 <= _1051;
        else
            _1052 <= _1049;
    end
    assign _1081 = _1052 & _1080;
    assign _1082 = _129 & _1081;
    assign write_enable_58 = _1082 & PHASE_13;
    assign _1087 = write_enable_58 | read_enable_48;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_28
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1087), .regcea(vdd), .wea(write_enable_58), .addra(address_58), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_49), .regceb(vdd), .web(write_enable_49), .addrb(address_49), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1094[131:131]), .sbiterrb(_1094[130:130]), .doutb(_1094[129:66]), .dbiterra(_1094[65:65]), .sbiterra(_1094[64:64]), .douta(_1094[63:0]) );
    assign _1095 = _1094[63:0];
    assign _1025 = ~ PHASE_13;
    assign _39 = _1025;
    always @(posedge _84) begin
        if (_82)
            PHASE_13 <= _1023;
        else
            if (_72)
                PHASE_13 <= _39;
    end
    assign _1107 = PHASE_13 ? _1106 : _1095;
    assign address_59 = _1280 ? _199 : _1275;
    assign write_enable_59 = _1273 & _1280;
    assign address_60 = _1280 ? _164 : _68;
    assign _1282 = ~ _1280;
    assign read_enable_49 = _1268 & _1282;
    assign _1280 = ~ PHASE_16;
    assign write_enable_60 = _1266 & _1280;
    assign _1284 = write_enable_60 | read_enable_49;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_29
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1284), .regcea(vdd), .wea(write_enable_60), .addra(address_60), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_59), .regceb(vdd), .web(write_enable_59), .addrb(address_59), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1289[131:131]), .sbiterrb(_1289[130:130]), .doutb(_1289[129:66]), .dbiterra(_1289[65:65]), .sbiterra(_1289[64:64]), .douta(_1289[63:0]) );
    assign _1290 = _1289[63:0];
    assign address_61 = PHASE_16 ? _199 : _1275;
    assign _1273 = _129 & _1236;
    assign write_enable_61 = _1273 & PHASE_16;
    assign _1198 = _1190[129:66];
    assign _1197 = _1177[129:66];
    assign _1199 = PHASE_14 ? _1198 : _1197;
    assign _1195 = _1147[129:66];
    assign _1194 = _1133[129:66];
    assign q1_4 = PHASE_15 ? _1195 : _1194;
    assign _1200 = _1114 ? _1199 : q1_4;
    assign address_62 = _1179 ? _1173 : _1172;
    assign _1185 = ~ _1179;
    assign read_enable_50 = _102 & _1185;
    assign address_63 = _1179 ? _60 : _1161;
    assign _1181 = ~ _1179;
    assign read_enable_51 = _102 & _1181;
    assign _1179 = ~ PHASE_14;
    assign write_enable_63 = _1150 & _1179;
    assign _1183 = write_enable_63 | read_enable_51;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_30
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1183), .regcea(vdd), .wea(write_enable_63), .addra(address_63), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_50), .regceb(vdd), .web(write_enable_62), .addrb(address_62), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1190[131:131]), .sbiterrb(_1190[130:130]), .doutb(_1190[129:66]), .dbiterra(_1190[65:65]), .sbiterra(_1190[64:64]), .douta(_1190[63:0]) );
    assign _1191 = _1190[63:0];
    assign _1171 = _172[5:5];
    assign _1170 = _172[4:4];
    assign _1169 = _172[3:3];
    assign _1168 = _172[2:2];
    assign _1167 = _172[1:1];
    assign _1166 = _172[0:0];
    assign _1172 = { _1166, _1167, _1168, _1169, _1170, _1171 };
    assign address_64 = PHASE_14 ? _1173 : _1172;
    assign _1163 = ~ PHASE_14;
    assign read_enable_52 = _102 & _1163;
    assign data_61 = wr_d2;
    assign _1160 = _137[5:5];
    assign _1159 = _137[4:4];
    assign _1158 = _137[3:3];
    assign _1157 = _137[2:2];
    assign _1156 = _137[1:1];
    assign _1155 = _137[0:0];
    assign _1161 = { _1155, _1156, _1157, _1158, _1159, _1160 };
    assign address_65 = PHASE_14 ? _60 : _1161;
    assign _1152 = ~ PHASE_14;
    assign read_enable_53 = _102 & _1152;
    assign _1150 = _62[2:2];
    assign write_enable_65 = _1150 & PHASE_14;
    assign _1154 = write_enable_65 | read_enable_53;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_31
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1154), .regcea(vdd), .wea(write_enable_65), .addra(address_65), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_52), .regceb(vdd), .web(write_enable_64), .addrb(address_64), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1177[131:131]), .sbiterrb(_1177[130:130]), .doutb(_1177[129:66]), .dbiterra(_1177[65:65]), .sbiterra(_1177[64:64]), .douta(_1177[63:0]) );
    assign _1178 = _1177[63:0];
    assign _1111 = ~ PHASE_14;
    assign _43 = _1111;
    always @(posedge _84) begin
        if (_82)
            PHASE_14 <= _1109;
        else
            if (_72)
                PHASE_14 <= _43;
    end
    assign _1192 = PHASE_14 ? _1191 : _1178;
    assign address_66 = _1135 ? _199 : _172;
    assign _1142 = ~ _1135;
    assign read_enable_54 = _102 & _1142;
    assign write_enable_66 = _1126 & _1135;
    assign _1144 = write_enable_66 | read_enable_54;
    assign address_67 = _1135 ? _164 : _137;
    assign _1137 = ~ _1135;
    assign read_enable_55 = _102 & _1137;
    assign _1135 = ~ PHASE_15;
    assign write_enable_67 = _1119 & _1135;
    assign _1139 = write_enable_67 | read_enable_55;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_32
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1139), .regcea(vdd), .wea(write_enable_67), .addra(address_67), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1144), .regceb(vdd), .web(write_enable_66), .addrb(address_66), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1147[131:131]), .sbiterrb(_1147[130:130]), .doutb(_1147[129:66]), .dbiterra(_1147[65:65]), .sbiterra(_1147[64:64]), .douta(_1147[63:0]) );
    assign _1148 = _1147[63:0];
    assign _1203 = _1202[127:64];
    assign data_63 = _1203;
    assign address_68 = PHASE_15 ? _199 : _172;
    assign _1128 = ~ PHASE_15;
    assign read_enable_56 = _102 & _1128;
    assign _1125 = ~ _130;
    assign _1126 = _129 & _1125;
    assign write_enable_68 = _1126 & PHASE_15;
    assign _1130 = write_enable_68 | read_enable_56;
    assign address_69 = PHASE_15 ? _164 : _137;
    assign _1121 = ~ PHASE_15;
    assign read_enable_57 = _102 & _1121;
    assign _1118 = ~ _130;
    assign _1119 = _129 & _1118;
    assign write_enable_69 = _1119 & PHASE_15;
    assign _1123 = write_enable_69 | read_enable_57;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_33
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1123), .regcea(vdd), .wea(write_enable_69), .addra(address_69), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1130), .regceb(vdd), .web(write_enable_68), .addrb(address_68), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1133[131:131]), .sbiterrb(_1133[130:130]), .doutb(_1133[129:66]), .dbiterra(_1133[65:65]), .sbiterra(_1133[64:64]), .douta(_1133[63:0]) );
    assign _1134 = _1133[63:0];
    assign _1204 = ~ PHASE_15;
    assign _45 = _1204;
    always @(posedge _84) begin
        if (_82)
            PHASE_15 <= _1116;
        else
            if (_99)
                PHASE_15 <= _45;
    end
    assign q0_4 = PHASE_15 ? _1148 : _1134;
    always @(posedge _84) begin
        if (_82)
            _1114 <= _1113;
        else
            _1114 <= _92;
    end
    assign _1193 = _1114 ? _1192 : q0_4;
    dp_1
        dp_1
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1193), .d2(_1200), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_1202[191:128]), .q2(_1202[127:64]), .q1(_1202[63:0]) );
    assign _1205 = _1202[63:0];
    assign data_67 = _1205;
    assign address_70 = PHASE_16 ? _164 : _68;
    assign _1269 = ~ PHASE_16;
    assign _1268 = _70[2:2];
    assign read_enable_58 = _1268 & _1269;
    always @(posedge _84) begin
        if (_82)
            _1239 <= _1238;
        else
            _1239 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _1242 <= _1241;
        else
            _1242 <= _1239;
    end
    always @(posedge _84) begin
        if (_82)
            _1245 <= _1244;
        else
            _1245 <= _1242;
    end
    always @(posedge _84) begin
        if (_82)
            _1248 <= _1247;
        else
            _1248 <= _1245;
    end
    always @(posedge _84) begin
        if (_82)
            _1251 <= _1250;
        else
            _1251 <= _1248;
    end
    always @(posedge _84) begin
        if (_82)
            _1254 <= _1253;
        else
            _1254 <= _1251;
    end
    always @(posedge _84) begin
        if (_82)
            _1257 <= _1256;
        else
            _1257 <= _1254;
    end
    always @(posedge _84) begin
        if (_82)
            _1260 <= _1259;
        else
            _1260 <= _1257;
    end
    always @(posedge _84) begin
        if (_82)
            _1263 <= _1262;
        else
            _1263 <= _1260;
    end
    assign _1264 = ~ _1263;
    always @(posedge _84) begin
        if (_82)
            _1212 <= _1211;
        else
            _1212 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1215 <= _1214;
        else
            _1215 <= _1212;
    end
    always @(posedge _84) begin
        if (_82)
            _1218 <= _1217;
        else
            _1218 <= _1215;
    end
    always @(posedge _84) begin
        if (_82)
            _1221 <= _1220;
        else
            _1221 <= _1218;
    end
    always @(posedge _84) begin
        if (_82)
            _1224 <= _1223;
        else
            _1224 <= _1221;
    end
    always @(posedge _84) begin
        if (_82)
            _1227 <= _1226;
        else
            _1227 <= _1224;
    end
    always @(posedge _84) begin
        if (_82)
            _1230 <= _1229;
        else
            _1230 <= _1227;
    end
    always @(posedge _84) begin
        if (_82)
            _1233 <= _1232;
        else
            _1233 <= _1230;
    end
    always @(posedge _84) begin
        if (_82)
            _1236 <= _1235;
        else
            _1236 <= _1233;
    end
    assign _1265 = _1236 & _1264;
    assign _1266 = _129 & _1265;
    assign write_enable_70 = _1266 & PHASE_16;
    assign _1271 = write_enable_70 | read_enable_58;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_34
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1271), .regcea(vdd), .wea(write_enable_70), .addra(address_70), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_61), .regceb(vdd), .web(write_enable_61), .addrb(address_61), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1278[131:131]), .sbiterrb(_1278[130:130]), .doutb(_1278[129:66]), .dbiterra(_1278[65:65]), .sbiterra(_1278[64:64]), .douta(_1278[63:0]) );
    assign _1279 = _1278[63:0];
    assign _1209 = ~ PHASE_16;
    assign _47 = _1209;
    always @(posedge _84) begin
        if (_82)
            PHASE_16 <= _1207;
        else
            if (_72)
                PHASE_16 <= _47;
    end
    assign _1291 = PHASE_16 ? _1290 : _1279;
    assign address_71 = _1464 ? _199 : _1459;
    assign write_enable_71 = _1457 & _1464;
    assign address_72 = _1464 ? _164 : _68;
    assign _1466 = ~ _1464;
    assign read_enable_59 = _1452 & _1466;
    assign _1464 = ~ PHASE_19;
    assign write_enable_72 = _1450 & _1464;
    assign _1468 = write_enable_72 | read_enable_59;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_35
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1468), .regcea(vdd), .wea(write_enable_72), .addra(address_72), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_71), .regceb(vdd), .web(write_enable_71), .addrb(address_71), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1473[131:131]), .sbiterrb(_1473[130:130]), .doutb(_1473[129:66]), .dbiterra(_1473[65:65]), .sbiterra(_1473[64:64]), .douta(_1473[63:0]) );
    assign _1474 = _1473[63:0];
    assign address_73 = PHASE_19 ? _199 : _1459;
    assign _1457 = _129 & _1420;
    assign write_enable_73 = _1457 & PHASE_19;
    assign _1382 = _1374[129:66];
    assign _1381 = _1361[129:66];
    assign _1383 = PHASE_17 ? _1382 : _1381;
    assign _1379 = _1331[129:66];
    assign _1378 = _1317[129:66];
    assign q1_5 = PHASE_18 ? _1379 : _1378;
    assign _1384 = _1298 ? _1383 : q1_5;
    assign address_74 = _1363 ? _1357 : _1356;
    assign _1369 = ~ _1363;
    assign read_enable_60 = _102 & _1369;
    assign address_75 = _1363 ? _60 : _1345;
    assign _1365 = ~ _1363;
    assign read_enable_61 = _102 & _1365;
    assign _1363 = ~ PHASE_17;
    assign write_enable_75 = _1334 & _1363;
    assign _1367 = write_enable_75 | read_enable_61;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_36
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1367), .regcea(vdd), .wea(write_enable_75), .addra(address_75), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_60), .regceb(vdd), .web(write_enable_74), .addrb(address_74), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1374[131:131]), .sbiterrb(_1374[130:130]), .doutb(_1374[129:66]), .dbiterra(_1374[65:65]), .sbiterra(_1374[64:64]), .douta(_1374[63:0]) );
    assign _1375 = _1374[63:0];
    assign _1355 = _172[5:5];
    assign _1354 = _172[4:4];
    assign _1353 = _172[3:3];
    assign _1352 = _172[2:2];
    assign _1351 = _172[1:1];
    assign _1350 = _172[0:0];
    assign _1356 = { _1350, _1351, _1352, _1353, _1354, _1355 };
    assign address_76 = PHASE_17 ? _1357 : _1356;
    assign _1347 = ~ PHASE_17;
    assign read_enable_62 = _102 & _1347;
    assign data_73 = wr_d1;
    assign _1344 = _137[5:5];
    assign _1343 = _137[4:4];
    assign _1342 = _137[3:3];
    assign _1341 = _137[2:2];
    assign _1340 = _137[1:1];
    assign _1339 = _137[0:0];
    assign _1345 = { _1339, _1340, _1341, _1342, _1343, _1344 };
    assign address_77 = PHASE_17 ? _60 : _1345;
    assign _1336 = ~ PHASE_17;
    assign read_enable_63 = _102 & _1336;
    assign _1334 = _62[1:1];
    assign write_enable_77 = _1334 & PHASE_17;
    assign _1338 = write_enable_77 | read_enable_63;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_37
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1338), .regcea(vdd), .wea(write_enable_77), .addra(address_77), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_62), .regceb(vdd), .web(write_enable_76), .addrb(address_76), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1361[131:131]), .sbiterrb(_1361[130:130]), .doutb(_1361[129:66]), .dbiterra(_1361[65:65]), .sbiterra(_1361[64:64]), .douta(_1361[63:0]) );
    assign _1362 = _1361[63:0];
    assign _1295 = ~ PHASE_17;
    assign _51 = _1295;
    always @(posedge _84) begin
        if (_82)
            PHASE_17 <= _1293;
        else
            if (_72)
                PHASE_17 <= _51;
    end
    assign _1376 = PHASE_17 ? _1375 : _1362;
    assign address_78 = _1319 ? _199 : _172;
    assign _1326 = ~ _1319;
    assign read_enable_64 = _102 & _1326;
    assign write_enable_78 = _1310 & _1319;
    assign _1328 = write_enable_78 | read_enable_64;
    assign address_79 = _1319 ? _164 : _137;
    assign _1321 = ~ _1319;
    assign read_enable_65 = _102 & _1321;
    assign _1319 = ~ PHASE_18;
    assign write_enable_79 = _1303 & _1319;
    assign _1323 = write_enable_79 | read_enable_65;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_38
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1323), .regcea(vdd), .wea(write_enable_79), .addra(address_79), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1328), .regceb(vdd), .web(write_enable_78), .addrb(address_78), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1331[131:131]), .sbiterrb(_1331[130:130]), .doutb(_1331[129:66]), .dbiterra(_1331[65:65]), .sbiterra(_1331[64:64]), .douta(_1331[63:0]) );
    assign _1332 = _1331[63:0];
    assign _1387 = _1386[127:64];
    assign data_75 = _1387;
    assign address_80 = PHASE_18 ? _199 : _172;
    assign _1312 = ~ PHASE_18;
    assign read_enable_66 = _102 & _1312;
    assign _1309 = ~ _130;
    assign _1310 = _129 & _1309;
    assign write_enable_80 = _1310 & PHASE_18;
    assign _1314 = write_enable_80 | read_enable_66;
    assign address_81 = PHASE_18 ? _164 : _137;
    assign _1305 = ~ PHASE_18;
    assign read_enable_67 = _102 & _1305;
    assign _1302 = ~ _130;
    assign _1303 = _129 & _1302;
    assign write_enable_81 = _1303 & PHASE_18;
    assign _1307 = write_enable_81 | read_enable_67;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_39
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1307), .regcea(vdd), .wea(write_enable_81), .addra(address_81), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1314), .regceb(vdd), .web(write_enable_80), .addrb(address_80), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1317[131:131]), .sbiterrb(_1317[130:130]), .doutb(_1317[129:66]), .dbiterra(_1317[65:65]), .sbiterra(_1317[64:64]), .douta(_1317[63:0]) );
    assign _1318 = _1317[63:0];
    assign _1388 = ~ PHASE_18;
    assign _53 = _1388;
    always @(posedge _84) begin
        if (_82)
            PHASE_18 <= _1300;
        else
            if (_99)
                PHASE_18 <= _53;
    end
    assign q0_5 = PHASE_18 ? _1332 : _1318;
    always @(posedge _84) begin
        if (_82)
            _1298 <= _1297;
        else
            _1298 <= _92;
    end
    assign _1377 = _1298 ? _1376 : q0_5;
    dp_0
        dp_0
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1377), .d2(_1384), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_1386[191:128]), .q2(_1386[127:64]), .q1(_1386[63:0]) );
    assign _1389 = _1386[63:0];
    assign data_79 = _1389;
    assign address_82 = PHASE_19 ? _164 : _68;
    assign _1453 = ~ PHASE_19;
    assign _1452 = _70[1:1];
    assign read_enable_68 = _1452 & _1453;
    always @(posedge _84) begin
        if (_82)
            _1423 <= _1422;
        else
            _1423 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _1426 <= _1425;
        else
            _1426 <= _1423;
    end
    always @(posedge _84) begin
        if (_82)
            _1429 <= _1428;
        else
            _1429 <= _1426;
    end
    always @(posedge _84) begin
        if (_82)
            _1432 <= _1431;
        else
            _1432 <= _1429;
    end
    always @(posedge _84) begin
        if (_82)
            _1435 <= _1434;
        else
            _1435 <= _1432;
    end
    always @(posedge _84) begin
        if (_82)
            _1438 <= _1437;
        else
            _1438 <= _1435;
    end
    always @(posedge _84) begin
        if (_82)
            _1441 <= _1440;
        else
            _1441 <= _1438;
    end
    always @(posedge _84) begin
        if (_82)
            _1444 <= _1443;
        else
            _1444 <= _1441;
    end
    always @(posedge _84) begin
        if (_82)
            _1447 <= _1446;
        else
            _1447 <= _1444;
    end
    assign _1448 = ~ _1447;
    always @(posedge _84) begin
        if (_82)
            _1396 <= _1395;
        else
            _1396 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1399 <= _1398;
        else
            _1399 <= _1396;
    end
    always @(posedge _84) begin
        if (_82)
            _1402 <= _1401;
        else
            _1402 <= _1399;
    end
    always @(posedge _84) begin
        if (_82)
            _1405 <= _1404;
        else
            _1405 <= _1402;
    end
    always @(posedge _84) begin
        if (_82)
            _1408 <= _1407;
        else
            _1408 <= _1405;
    end
    always @(posedge _84) begin
        if (_82)
            _1411 <= _1410;
        else
            _1411 <= _1408;
    end
    always @(posedge _84) begin
        if (_82)
            _1414 <= _1413;
        else
            _1414 <= _1411;
    end
    always @(posedge _84) begin
        if (_82)
            _1417 <= _1416;
        else
            _1417 <= _1414;
    end
    always @(posedge _84) begin
        if (_82)
            _1420 <= _1419;
        else
            _1420 <= _1417;
    end
    assign _1449 = _1420 & _1448;
    assign _1450 = _129 & _1449;
    assign write_enable_82 = _1450 & PHASE_19;
    assign _1455 = write_enable_82 | read_enable_68;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_40
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1455), .regcea(vdd), .wea(write_enable_82), .addra(address_82), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_73), .regceb(vdd), .web(write_enable_73), .addrb(address_73), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1462[131:131]), .sbiterrb(_1462[130:130]), .doutb(_1462[129:66]), .dbiterra(_1462[65:65]), .sbiterra(_1462[64:64]), .douta(_1462[63:0]) );
    assign _1463 = _1462[63:0];
    assign _1393 = ~ PHASE_19;
    assign _55 = _1393;
    always @(posedge _84) begin
        if (_82)
            PHASE_19 <= _1391;
        else
            if (_72)
                PHASE_19 <= _55;
    end
    assign _1475 = PHASE_19 ? _1474 : _1463;
    assign address_83 = _1648 ? _199 : _1643;
    assign write_enable_83 = _1641 & _1648;
    assign address_84 = _1648 ? _164 : _68;
    assign _1650 = ~ _1648;
    assign read_enable_69 = _1636 & _1650;
    assign _1648 = ~ PHASE_22;
    assign write_enable_84 = _1634 & _1648;
    assign _1652 = write_enable_84 | read_enable_69;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_41
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1652), .regcea(vdd), .wea(write_enable_84), .addra(address_84), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_83), .regceb(vdd), .web(write_enable_83), .addrb(address_83), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1657[131:131]), .sbiterrb(_1657[130:130]), .doutb(_1657[129:66]), .dbiterra(_1657[65:65]), .sbiterra(_1657[64:64]), .douta(_1657[63:0]) );
    assign _1658 = _1657[63:0];
    assign address_85 = PHASE_22 ? _199 : _1643;
    assign _1641 = _129 & _1604;
    assign write_enable_85 = _1641 & PHASE_22;
    assign _280 = _91[490:487];
    assign _279 = _91[486:486];
    assign _277 = _91[482:482];
    assign _276 = _91[481:418];
    assign _275 = _91[417:354];
    assign _274 = _91[353:290];
    assign _273 = _91[289:226];
    assign _272 = _91[225:162];
    assign _271 = _91[161:98];
    assign _270 = _91[97:34];
    assign _1566 = _1558[129:66];
    assign _1565 = _1545[129:66];
    assign _1567 = PHASE_20 ? _1566 : _1565;
    assign _1563 = _1515[129:66];
    assign _1562 = _1501[129:66];
    assign q1_6 = PHASE_21 ? _1563 : _1562;
    assign _1568 = _1482 ? _1567 : q1_6;
    assign address_86 = _1547 ? _1541 : _1540;
    assign _1553 = ~ _1547;
    assign read_enable_70 = _102 & _1553;
    assign address_87 = _1547 ? _60 : _1529;
    assign _1549 = ~ _1547;
    assign read_enable_71 = _102 & _1549;
    assign _1547 = ~ PHASE_20;
    assign write_enable_87 = _1518 & _1547;
    assign _1551 = write_enable_87 | read_enable_71;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_42
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1551), .regcea(vdd), .wea(write_enable_87), .addra(address_87), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_70), .regceb(vdd), .web(write_enable_86), .addrb(address_86), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1558[131:131]), .sbiterrb(_1558[130:130]), .doutb(_1558[129:66]), .dbiterra(_1558[65:65]), .sbiterra(_1558[64:64]), .douta(_1558[63:0]) );
    assign _1559 = _1558[63:0];
    assign _1539 = _172[5:5];
    assign _1538 = _172[4:4];
    assign _1537 = _172[3:3];
    assign _1536 = _172[2:2];
    assign _1535 = _172[1:1];
    assign _1534 = _172[0:0];
    assign _1540 = { _1534, _1535, _1536, _1537, _1538, _1539 };
    assign address_88 = PHASE_20 ? _1541 : _1540;
    assign _1531 = ~ PHASE_20;
    assign read_enable_72 = _102 & _1531;
    assign data_85 = wr_d0;
    assign _60 = wr_addr;
    assign _1528 = _137[5:5];
    assign _1527 = _137[4:4];
    assign _1526 = _137[3:3];
    assign _1525 = _137[2:2];
    assign _1524 = _137[1:1];
    assign _1523 = _137[0:0];
    assign _1529 = { _1523, _1524, _1525, _1526, _1527, _1528 };
    assign address_89 = PHASE_20 ? _60 : _1529;
    assign _1520 = ~ PHASE_20;
    assign read_enable_73 = _102 & _1520;
    assign _62 = wr_en;
    assign _1518 = _62[0:0];
    assign write_enable_89 = _1518 & PHASE_20;
    assign _1522 = write_enable_89 | read_enable_73;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_43
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1522), .regcea(vdd), .wea(write_enable_89), .addra(address_89), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_72), .regceb(vdd), .web(write_enable_88), .addrb(address_88), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1545[131:131]), .sbiterrb(_1545[130:130]), .doutb(_1545[129:66]), .dbiterra(_1545[65:65]), .sbiterra(_1545[64:64]), .douta(_1545[63:0]) );
    assign _1546 = _1545[63:0];
    assign _1479 = ~ PHASE_20;
    assign _63 = _1479;
    always @(posedge _84) begin
        if (_82)
            PHASE_20 <= _1477;
        else
            if (_72)
                PHASE_20 <= _63;
    end
    assign _1560 = PHASE_20 ? _1559 : _1546;
    assign address_90 = _1503 ? _199 : _172;
    assign _1510 = ~ _1503;
    assign read_enable_74 = _102 & _1510;
    assign write_enable_90 = _1494 & _1503;
    assign _1512 = write_enable_90 | read_enable_74;
    assign address_91 = _1503 ? _164 : _137;
    assign _1505 = ~ _1503;
    assign read_enable_75 = _102 & _1505;
    assign _1503 = ~ PHASE_21;
    assign write_enable_91 = _1487 & _1503;
    assign _1507 = write_enable_91 | read_enable_75;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_44
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1507), .regcea(vdd), .wea(write_enable_91), .addra(address_91), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1512), .regceb(vdd), .web(write_enable_90), .addrb(address_90), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1515[131:131]), .sbiterrb(_1515[130:130]), .doutb(_1515[129:66]), .dbiterra(_1515[65:65]), .sbiterra(_1515[64:64]), .douta(_1515[63:0]) );
    assign _1516 = _1515[63:0];
    assign _1571 = _1570[127:64];
    assign data_87 = _1571;
    always @(posedge _84) begin
        if (_82)
            _175 <= _174;
        else
            _175 <= _172;
    end
    always @(posedge _84) begin
        if (_82)
            _178 <= _177;
        else
            _178 <= _175;
    end
    always @(posedge _84) begin
        if (_82)
            _181 <= _180;
        else
            _181 <= _178;
    end
    always @(posedge _84) begin
        if (_82)
            _184 <= _183;
        else
            _184 <= _181;
    end
    always @(posedge _84) begin
        if (_82)
            _187 <= _186;
        else
            _187 <= _184;
    end
    always @(posedge _84) begin
        if (_82)
            _190 <= _189;
        else
            _190 <= _187;
    end
    always @(posedge _84) begin
        if (_82)
            _193 <= _192;
        else
            _193 <= _190;
    end
    always @(posedge _84) begin
        if (_82)
            _196 <= _195;
        else
            _196 <= _193;
    end
    always @(posedge _84) begin
        if (_82)
            _199 <= _198;
        else
            _199 <= _196;
    end
    assign _172 = _91[33:28];
    assign address_92 = PHASE_21 ? _199 : _172;
    assign _1496 = ~ PHASE_21;
    assign read_enable_76 = _102 & _1496;
    assign _1493 = ~ _130;
    assign _1494 = _129 & _1493;
    assign write_enable_92 = _1494 & PHASE_21;
    assign _1498 = write_enable_92 | read_enable_76;
    assign address_93 = PHASE_21 ? _164 : _137;
    assign _1489 = ~ PHASE_21;
    assign read_enable_77 = _102 & _1489;
    assign _1486 = ~ _130;
    assign _1487 = _129 & _1486;
    assign write_enable_93 = _1487 & PHASE_21;
    assign _1491 = write_enable_93 | read_enable_77;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_45
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1491), .regcea(vdd), .wea(write_enable_93), .addra(address_93), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1498), .regceb(vdd), .web(write_enable_92), .addrb(address_92), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1501[131:131]), .sbiterrb(_1501[130:130]), .doutb(_1501[129:66]), .dbiterra(_1501[65:65]), .sbiterra(_1501[64:64]), .douta(_1501[63:0]) );
    assign _1502 = _1501[63:0];
    assign _99 = _91[492:492];
    assign _1572 = ~ PHASE_21;
    assign _65 = _1572;
    always @(posedge _84) begin
        if (_82)
            PHASE_21 <= _1484;
        else
            if (_99)
                PHASE_21 <= _65;
    end
    assign q0_6 = PHASE_21 ? _1516 : _1502;
    assign _92 = _91[483:483];
    always @(posedge _84) begin
        if (_82)
            _1482 <= _1481;
        else
            _1482 <= _92;
    end
    assign _1561 = _1482 ? _1560 : q0_6;
    dp
        dp
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1561), .d2(_1568), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_1570[191:128]), .q2(_1570[127:64]), .q1(_1570[63:0]) );
    assign _1573 = _1570[63:0];
    assign data_91 = _1573;
    assign _137 = _91[27:22];
    always @(posedge _84) begin
        if (_82)
            _140 <= _139;
        else
            _140 <= _137;
    end
    always @(posedge _84) begin
        if (_82)
            _143 <= _142;
        else
            _143 <= _140;
    end
    always @(posedge _84) begin
        if (_82)
            _146 <= _145;
        else
            _146 <= _143;
    end
    always @(posedge _84) begin
        if (_82)
            _149 <= _148;
        else
            _149 <= _146;
    end
    always @(posedge _84) begin
        if (_82)
            _152 <= _151;
        else
            _152 <= _149;
    end
    always @(posedge _84) begin
        if (_82)
            _155 <= _154;
        else
            _155 <= _152;
    end
    always @(posedge _84) begin
        if (_82)
            _158 <= _157;
        else
            _158 <= _155;
    end
    always @(posedge _84) begin
        if (_82)
            _161 <= _160;
        else
            _161 <= _158;
    end
    always @(posedge _84) begin
        if (_82)
            _164 <= _163;
        else
            _164 <= _161;
    end
    assign _68 = rd_addr;
    assign address_94 = PHASE_22 ? _164 : _68;
    assign _1637 = ~ PHASE_22;
    assign _70 = rd_en;
    assign _1636 = _70[0:0];
    assign read_enable_78 = _1636 & _1637;
    assign _278 = _91[485:485];
    always @(posedge _84) begin
        if (_82)
            _1607 <= _1606;
        else
            _1607 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _1610 <= _1609;
        else
            _1610 <= _1607;
    end
    always @(posedge _84) begin
        if (_82)
            _1613 <= _1612;
        else
            _1613 <= _1610;
    end
    always @(posedge _84) begin
        if (_82)
            _1616 <= _1615;
        else
            _1616 <= _1613;
    end
    always @(posedge _84) begin
        if (_82)
            _1619 <= _1618;
        else
            _1619 <= _1616;
    end
    always @(posedge _84) begin
        if (_82)
            _1622 <= _1621;
        else
            _1622 <= _1619;
    end
    always @(posedge _84) begin
        if (_82)
            _1625 <= _1624;
        else
            _1625 <= _1622;
    end
    always @(posedge _84) begin
        if (_82)
            _1628 <= _1627;
        else
            _1628 <= _1625;
    end
    always @(posedge _84) begin
        if (_82)
            _1631 <= _1630;
        else
            _1631 <= _1628;
    end
    assign _1632 = ~ _1631;
    assign _130 = _91[484:484];
    always @(posedge _84) begin
        if (_82)
            _1580 <= _1579;
        else
            _1580 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1583 <= _1582;
        else
            _1583 <= _1580;
    end
    always @(posedge _84) begin
        if (_82)
            _1586 <= _1585;
        else
            _1586 <= _1583;
    end
    always @(posedge _84) begin
        if (_82)
            _1589 <= _1588;
        else
            _1589 <= _1586;
    end
    always @(posedge _84) begin
        if (_82)
            _1592 <= _1591;
        else
            _1592 <= _1589;
    end
    always @(posedge _84) begin
        if (_82)
            _1595 <= _1594;
        else
            _1595 <= _1592;
    end
    always @(posedge _84) begin
        if (_82)
            _1598 <= _1597;
        else
            _1598 <= _1595;
    end
    always @(posedge _84) begin
        if (_82)
            _1601 <= _1600;
        else
            _1601 <= _1598;
    end
    always @(posedge _84) begin
        if (_82)
            _1604 <= _1603;
        else
            _1604 <= _1601;
    end
    assign _1633 = _1604 & _1632;
    assign _102 = _91[491:491];
    always @(posedge _84) begin
        if (_82)
            _105 <= _104;
        else
            _105 <= _102;
    end
    always @(posedge _84) begin
        if (_82)
            _108 <= _107;
        else
            _108 <= _105;
    end
    always @(posedge _84) begin
        if (_82)
            _111 <= _110;
        else
            _111 <= _108;
    end
    always @(posedge _84) begin
        if (_82)
            _114 <= _113;
        else
            _114 <= _111;
    end
    always @(posedge _84) begin
        if (_82)
            _117 <= _116;
        else
            _117 <= _114;
    end
    always @(posedge _84) begin
        if (_82)
            _120 <= _119;
        else
            _120 <= _117;
    end
    always @(posedge _84) begin
        if (_82)
            _123 <= _122;
        else
            _123 <= _120;
    end
    always @(posedge _84) begin
        if (_82)
            _126 <= _125;
        else
            _126 <= _123;
    end
    always @(posedge _84) begin
        if (_82)
            _129 <= _128;
        else
            _129 <= _126;
    end
    assign _1634 = _129 & _1633;
    assign write_enable_94 = _1634 & PHASE_22;
    assign _1639 = write_enable_94 | read_enable_78;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_46
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1639), .regcea(vdd), .wea(write_enable_94), .addra(address_94), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_85), .regceb(vdd), .web(write_enable_85), .addrb(address_85), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1646[131:131]), .sbiterrb(_1646[130:130]), .doutb(_1646[129:66]), .dbiterra(_1646[65:65]), .sbiterra(_1646[64:64]), .douta(_1646[63:0]) );
    assign _1647 = _1646[63:0];
    assign _72 = flip;
    assign _1577 = ~ PHASE_22;
    assign _73 = _1577;
    always @(posedge _84) begin
        if (_82)
            PHASE_22 <= _1575;
        else
            if (_72)
                PHASE_22 <= _73;
    end
    assign _1659 = PHASE_22 ? _1658 : _1647;
    assign _76 = first_4step_pass;
    assign _78 = first_iter;
    assign _80 = start;
    assign _82 = clear;
    assign _84 = clock;
    ctrl
        ctrl
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .first_4step_pass(_76), .flip(_91[492:492]), .read_write_enable(_91[491:491]), .index(_91[490:487]), .valid(_91[486:486]), .twiddle_stage(_91[485:485]), .last_stage(_91[484:484]), .first_stage(_91[483:483]), .start_twiddles(_91[482:482]), .omegas6(_91[481:418]), .omegas5(_91[417:354]), .omegas4(_91[353:290]), .omegas3(_91[289:226]), .omegas2(_91[225:162]), .omegas1(_91[161:98]), .omegas0(_91[97:34]), .addr2(_91[33:28]), .addr1(_91[27:22]), .m(_91[21:16]), .k(_91[15:10]), .j(_91[9:4]), .i(_91[3:1]), .done_(_91[0:0]) );
    assign _1660 = _91[0:0];

    /* aliases */
    assign data_0 = data;
    assign data_2 = data_1;
    assign data_4 = data_3;
    assign data_5 = data_3;
    assign data_6 = data_3;
    assign data_8 = data_7;
    assign data_9 = data_7;
    assign data_10 = data_7;
    assign data_12 = data_11;
    assign data_14 = data_13;
    assign data_16 = data_15;
    assign data_17 = data_15;
    assign data_18 = data_15;
    assign data_20 = data_19;
    assign data_21 = data_19;
    assign data_22 = data_19;
    assign data_24 = data_23;
    assign data_26 = data_25;
    assign data_28 = data_27;
    assign data_29 = data_27;
    assign data_30 = data_27;
    assign data_32 = data_31;
    assign data_33 = data_31;
    assign data_34 = data_31;
    assign data_36 = data_35;
    assign data_38 = data_37;
    assign data_40 = data_39;
    assign data_41 = data_39;
    assign data_42 = data_39;
    assign data_44 = data_43;
    assign data_45 = data_43;
    assign data_46 = data_43;
    assign data_48 = data_47;
    assign data_50 = data_49;
    assign data_52 = data_51;
    assign data_53 = data_51;
    assign data_54 = data_51;
    assign data_56 = data_55;
    assign data_57 = data_55;
    assign data_58 = data_55;
    assign data_60 = data_59;
    assign data_62 = data_61;
    assign data_64 = data_63;
    assign data_65 = data_63;
    assign data_66 = data_63;
    assign data_68 = data_67;
    assign data_69 = data_67;
    assign data_70 = data_67;
    assign data_72 = data_71;
    assign data_74 = data_73;
    assign data_76 = data_75;
    assign data_77 = data_75;
    assign data_78 = data_75;
    assign data_80 = data_79;
    assign data_81 = data_79;
    assign data_82 = data_79;
    assign data_84 = data_83;
    assign data_86 = data_85;
    assign data_88 = data_87;
    assign data_89 = data_87;
    assign data_90 = data_87;
    assign data_92 = data_91;
    assign data_93 = data_91;
    assign data_94 = data_91;

    /* output assignments */
    assign done_ = _1660;
    assign rd_q0 = _1659;
    assign rd_q1 = _1475;
    assign rd_q2 = _1291;
    assign rd_q3 = _1107;
    assign rd_q4 = _923;
    assign rd_q5 = _739;
    assign rd_q6 = _555;
    assign rd_q7 = _371;

endmodule
module dp_7 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1001010110000011011011011110011100001111001100011100101111111010;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0000001111101000110111111101001001001110100011100111100000011111;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1100100001000011111100010110001010010100011000001011010101010001;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1011101000100101111010110101110011010001100101110000101011101011;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1011111101111001000101000011110011100110000011001010100101100110;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0001100100000101110100000010101001011100010000010001111101001110;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_8 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0101011011000110011100011000111110000111111100001101111000100011;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0111010010100011111001001101111110000010101010011101010011011100;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1001101100100100010111100000100001010011101110110101011011001110;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1110010100001110110001011011010111010011000010010011010110000000;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0101001110100110001000001111011110000111100111011011010111100001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0011101010100111000001000000100000001000111011011010110011010101;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1001110001100110000010001101010010111100110001111111101000100100;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_9 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0101011011101100000111100011111011111011000001010000001000001010;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0011100110101111101011010110110000110010100010110001011011110110;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1111111101011100001000000110011010110000001001110010101101001011;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1100100001000011111100010110001010010100011000001011010101010001;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0000001101001101110010111010010110001010110001010000000000111110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0011110110100000010111111110111001110000110001001111001010111010;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0111101001011001000101011001010111100110011111000010011111101000;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_10 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1001001001111111110101011000110110001111101011011001001101000000;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1111101010111110101001111000110111010110001001011011111111101111;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0001101010101101011111100110110011000101010001110000001110101000;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0100101110110010101100100000100001100011101000000110001110100010;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0110001000001000100101110011100101100010001000000001101110100011;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1010111010000110001000110110000101111000100111001100001010010101;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1010001011011001011001000100001001100101001010111001000111100101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_11 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0011001010101001010101000011100000101111110100000000100010101001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1010001101110111101111000010110101111101000101111110101011000110;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0011100110101111101011010110110000110010100010110001011011110110;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0000001111101000110111111101001001001110100011100111100000011111;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1110010100001110110001011011010111010011000010010011010110000000;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1011101000100101111010110101110011010001100101110000101011101011;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0110000010000100111001101000010001011010100100010010111101001101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_12 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1010000111101011011011000100001100101100111011111000010000010011;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1010000011011100010101000100001100110010011011110100111011000101;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0011000010100111001001111100101010011110010101110011001010111100;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0101110010000010010001101000010101000000100001101011001000100011;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0111010100000000110110011100011001101010010111101111110100110001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0000011100001011110100010000110110100011110110100100101101101110;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0110010011100000101001001101100100011100010001000101101011010010;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_13 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1011001100010001110110111110110011110001011101001011011101111001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0011001010101001010101000011100000101111110100000000100010101001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0101011011101100000111100011111011111011000001010000001000001010;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1001010110000011011011011110011100001111001100011100101111111010;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0110110110111110101101111110000000100110100001110010111000111001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0101010011010111101011100001010011111111011110000011001100001001;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1110111110011011001000010110000110000111101001101001011101000111;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_14 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0100110101000101100110100100101010000010100001001110100110001011;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0111001100001110001111011101000101111010000101110111100100101011;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0000001001111011000100111011001010010011010011011101111001111100;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0011100110101111101011010110110000110010100010110001011011110110;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1001101100100100010111100000100001010011101110110101011011001110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0000001101001101110010111010010110001010110001010000000000111110;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1110000001000010100010111011011100101110110101110011010000101110;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module parallel_cores_0 (
    wr_d7,
    wr_d6,
    wr_d5,
    wr_d4,
    wr_d3,
    wr_d2,
    wr_d1,
    wr_d0,
    wr_addr,
    wr_en,
    rd_addr,
    rd_en,
    flip,
    first_4step_pass,
    first_iter,
    start,
    clear,
    clock,
    done_,
    rd_q0,
    rd_q1,
    rd_q2,
    rd_q3,
    rd_q4,
    rd_q5,
    rd_q6,
    rd_q7
);

    input [63:0] wr_d7;
    input [63:0] wr_d6;
    input [63:0] wr_d5;
    input [63:0] wr_d4;
    input [63:0] wr_d3;
    input [63:0] wr_d2;
    input [63:0] wr_d1;
    input [63:0] wr_d0;
    input [5:0] wr_addr;
    input [7:0] wr_en;
    input [5:0] rd_addr;
    input [7:0] rd_en;
    input flip;
    input first_4step_pass;
    input first_iter;
    input start;
    input clear;
    input clock;
    output done_;
    output [63:0] rd_q0;
    output [63:0] rd_q1;
    output [63:0] rd_q2;
    output [63:0] rd_q3;
    output [63:0] rd_q4;
    output [63:0] rd_q5;
    output [63:0] rd_q6;
    output [63:0] rd_q7;

    /* signal declarations */
    wire [5:0] address;
    wire write_enable;
    wire [5:0] address_0;
    wire _362;
    wire read_enable;
    wire _360;
    wire write_enable_0;
    wire _364;
    wire [131:0] _369;
    wire [63:0] _370;
    wire [5:0] _355 = 6'b000000;
    wire [5:0] address_1;
    wire _353;
    wire write_enable_1;
    wire [63:0] _267;
    wire [63:0] _266;
    wire [63:0] _268;
    wire [63:0] _264;
    wire [63:0] _263;
    wire [63:0] q1;
    wire [63:0] _269;
    wire [5:0] address_2;
    wire write_enable_2 = 1'b0;
    wire _254;
    wire read_enable_0;
    wire [5:0] address_3;
    wire _250;
    wire read_enable_1;
    wire _248;
    wire write_enable_3;
    wire _252;
    wire [131:0] _259;
    wire [63:0] _260;
    wire [63:0] data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_0;
    wire [5:0] _242 = 6'b000000;
    wire _240;
    wire _239;
    wire _238;
    wire _237;
    wire _236;
    wire _235;
    wire [5:0] _241;
    wire [5:0] address_4;
    wire write_enable_4 = 1'b0;
    wire _232;
    wire read_enable_2;
    wire [63:0] data_1;
    wire [63:0] data_2;
    wire _229;
    wire _228;
    wire _227;
    wire _226;
    wire _225;
    wire _224;
    wire [5:0] _230;
    wire [5:0] address_5;
    wire _221;
    wire read_enable_3;
    wire _219;
    wire write_enable_5;
    wire _223;
    wire [131:0] _246;
    wire [63:0] _247;
    wire _87 = 1'b0;
    wire _86 = 1'b0;
    wire _89;
    wire _3;
    reg PHASE;
    wire [63:0] _261;
    wire [5:0] address_6;
    wire _211;
    wire read_enable_4;
    wire write_enable_6;
    wire _213;
    wire [5:0] address_7;
    wire _206;
    wire read_enable_5;
    wire _204;
    wire write_enable_7;
    wire _208;
    wire [131:0] _216;
    wire [63:0] _217;
    wire [63:0] _283;
    wire [63:0] data_3;
    wire [63:0] data_4;
    wire [63:0] data_5;
    wire [63:0] data_6;
    wire [5:0] address_8;
    wire _169;
    wire read_enable_6;
    wire _166;
    wire _167;
    wire write_enable_8;
    wire _171;
    wire [5:0] address_9;
    wire _134;
    wire read_enable_7;
    wire _131;
    wire _132;
    wire write_enable_9;
    wire _136;
    wire [131:0] _202;
    wire [63:0] _203;
    wire _98 = 1'b0;
    wire _97 = 1'b0;
    wire _284;
    wire _5;
    reg PHASE_0;
    wire [63:0] q0;
    wire _94 = 1'b0;
    wire _93 = 1'b0;
    reg _96;
    wire [63:0] _262;
    wire [191:0] _282;
    wire [63:0] _285;
    wire [63:0] data_7;
    wire [63:0] data_8;
    wire [63:0] data_9;
    wire [63:0] data_10;
    wire [5:0] address_10;
    wire _349;
    wire _348;
    wire read_enable_8;
    wire _342 = 1'b0;
    wire _341 = 1'b0;
    wire _339 = 1'b0;
    wire _338 = 1'b0;
    wire _336 = 1'b0;
    wire _335 = 1'b0;
    wire _333 = 1'b0;
    wire _332 = 1'b0;
    wire _330 = 1'b0;
    wire _329 = 1'b0;
    wire _327 = 1'b0;
    wire _326 = 1'b0;
    wire _324 = 1'b0;
    wire _323 = 1'b0;
    wire _321 = 1'b0;
    wire _320 = 1'b0;
    wire _318 = 1'b0;
    wire _317 = 1'b0;
    reg _319;
    reg _322;
    reg _325;
    reg _328;
    reg _331;
    reg _334;
    reg _337;
    reg _340;
    reg _343;
    wire _344;
    wire _315 = 1'b0;
    wire _314 = 1'b0;
    wire _312 = 1'b0;
    wire _311 = 1'b0;
    wire _309 = 1'b0;
    wire _308 = 1'b0;
    wire _306 = 1'b0;
    wire _305 = 1'b0;
    wire _303 = 1'b0;
    wire _302 = 1'b0;
    wire _300 = 1'b0;
    wire _299 = 1'b0;
    wire _297 = 1'b0;
    wire _296 = 1'b0;
    wire _294 = 1'b0;
    wire _293 = 1'b0;
    wire _291 = 1'b0;
    wire _290 = 1'b0;
    reg _292;
    reg _295;
    reg _298;
    reg _301;
    reg _304;
    reg _307;
    reg _310;
    reg _313;
    reg _316;
    wire _345;
    wire _346;
    wire write_enable_10;
    wire _351;
    wire [131:0] _358;
    wire [63:0] _359;
    wire _287 = 1'b0;
    wire _286 = 1'b0;
    wire _289;
    wire _7;
    reg PHASE_1;
    wire [63:0] _371;
    wire [5:0] address_11;
    wire write_enable_11;
    wire [5:0] address_12;
    wire _546;
    wire read_enable_9;
    wire _544;
    wire write_enable_12;
    wire _548;
    wire [131:0] _553;
    wire [63:0] _554;
    wire [5:0] _539 = 6'b000000;
    wire [5:0] address_13;
    wire _537;
    wire write_enable_13;
    wire [63:0] _462;
    wire [63:0] _461;
    wire [63:0] _463;
    wire [63:0] _459;
    wire [63:0] _458;
    wire [63:0] q1_0;
    wire [63:0] _464;
    wire [5:0] address_14;
    wire write_enable_14 = 1'b0;
    wire _449;
    wire read_enable_10;
    wire [5:0] address_15;
    wire _445;
    wire read_enable_11;
    wire _443;
    wire write_enable_15;
    wire _447;
    wire [131:0] _454;
    wire [63:0] _455;
    wire [63:0] data_11 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_12;
    wire [5:0] _437 = 6'b000000;
    wire _435;
    wire _434;
    wire _433;
    wire _432;
    wire _431;
    wire _430;
    wire [5:0] _436;
    wire [5:0] address_16;
    wire write_enable_16 = 1'b0;
    wire _427;
    wire read_enable_12;
    wire [63:0] data_13;
    wire [63:0] data_14;
    wire _424;
    wire _423;
    wire _422;
    wire _421;
    wire _420;
    wire _419;
    wire [5:0] _425;
    wire [5:0] address_17;
    wire _416;
    wire read_enable_13;
    wire _414;
    wire write_enable_17;
    wire _418;
    wire [131:0] _441;
    wire [63:0] _442;
    wire _373 = 1'b0;
    wire _372 = 1'b0;
    wire _375;
    wire _11;
    reg PHASE_2;
    wire [63:0] _456;
    wire [5:0] address_18;
    wire _406;
    wire read_enable_14;
    wire write_enable_18;
    wire _408;
    wire [5:0] address_19;
    wire _401;
    wire read_enable_15;
    wire _399;
    wire write_enable_19;
    wire _403;
    wire [131:0] _411;
    wire [63:0] _412;
    wire [63:0] _467;
    wire [63:0] data_15;
    wire [63:0] data_16;
    wire [63:0] data_17;
    wire [63:0] data_18;
    wire [5:0] address_20;
    wire _392;
    wire read_enable_16;
    wire _389;
    wire _390;
    wire write_enable_20;
    wire _394;
    wire [5:0] address_21;
    wire _385;
    wire read_enable_17;
    wire _382;
    wire _383;
    wire write_enable_21;
    wire _387;
    wire [131:0] _397;
    wire [63:0] _398;
    wire _380 = 1'b0;
    wire _379 = 1'b0;
    wire _468;
    wire _13;
    reg PHASE_3;
    wire [63:0] q0_0;
    wire _377 = 1'b0;
    wire _376 = 1'b0;
    reg _378;
    wire [63:0] _457;
    wire [191:0] _466;
    wire [63:0] _469;
    wire [63:0] data_19;
    wire [63:0] data_20;
    wire [63:0] data_21;
    wire [63:0] data_22;
    wire [5:0] address_22;
    wire _533;
    wire _532;
    wire read_enable_18;
    wire _526 = 1'b0;
    wire _525 = 1'b0;
    wire _523 = 1'b0;
    wire _522 = 1'b0;
    wire _520 = 1'b0;
    wire _519 = 1'b0;
    wire _517 = 1'b0;
    wire _516 = 1'b0;
    wire _514 = 1'b0;
    wire _513 = 1'b0;
    wire _511 = 1'b0;
    wire _510 = 1'b0;
    wire _508 = 1'b0;
    wire _507 = 1'b0;
    wire _505 = 1'b0;
    wire _504 = 1'b0;
    wire _502 = 1'b0;
    wire _501 = 1'b0;
    reg _503;
    reg _506;
    reg _509;
    reg _512;
    reg _515;
    reg _518;
    reg _521;
    reg _524;
    reg _527;
    wire _528;
    wire _499 = 1'b0;
    wire _498 = 1'b0;
    wire _496 = 1'b0;
    wire _495 = 1'b0;
    wire _493 = 1'b0;
    wire _492 = 1'b0;
    wire _490 = 1'b0;
    wire _489 = 1'b0;
    wire _487 = 1'b0;
    wire _486 = 1'b0;
    wire _484 = 1'b0;
    wire _483 = 1'b0;
    wire _481 = 1'b0;
    wire _480 = 1'b0;
    wire _478 = 1'b0;
    wire _477 = 1'b0;
    wire _475 = 1'b0;
    wire _474 = 1'b0;
    reg _476;
    reg _479;
    reg _482;
    reg _485;
    reg _488;
    reg _491;
    reg _494;
    reg _497;
    reg _500;
    wire _529;
    wire _530;
    wire write_enable_22;
    wire _535;
    wire [131:0] _542;
    wire [63:0] _543;
    wire _471 = 1'b0;
    wire _470 = 1'b0;
    wire _473;
    wire _15;
    reg PHASE_4;
    wire [63:0] _555;
    wire [5:0] address_23;
    wire write_enable_23;
    wire [5:0] address_24;
    wire _730;
    wire read_enable_19;
    wire _728;
    wire write_enable_24;
    wire _732;
    wire [131:0] _737;
    wire [63:0] _738;
    wire [5:0] _723 = 6'b000000;
    wire [5:0] address_25;
    wire _721;
    wire write_enable_25;
    wire [63:0] _646;
    wire [63:0] _645;
    wire [63:0] _647;
    wire [63:0] _643;
    wire [63:0] _642;
    wire [63:0] q1_1;
    wire [63:0] _648;
    wire [5:0] address_26;
    wire write_enable_26 = 1'b0;
    wire _633;
    wire read_enable_20;
    wire [5:0] address_27;
    wire _629;
    wire read_enable_21;
    wire _627;
    wire write_enable_27;
    wire _631;
    wire [131:0] _638;
    wire [63:0] _639;
    wire [63:0] data_23 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_24;
    wire [5:0] _621 = 6'b000000;
    wire _619;
    wire _618;
    wire _617;
    wire _616;
    wire _615;
    wire _614;
    wire [5:0] _620;
    wire [5:0] address_28;
    wire write_enable_28 = 1'b0;
    wire _611;
    wire read_enable_22;
    wire [63:0] data_25;
    wire [63:0] data_26;
    wire _608;
    wire _607;
    wire _606;
    wire _605;
    wire _604;
    wire _603;
    wire [5:0] _609;
    wire [5:0] address_29;
    wire _600;
    wire read_enable_23;
    wire _598;
    wire write_enable_29;
    wire _602;
    wire [131:0] _625;
    wire [63:0] _626;
    wire _557 = 1'b0;
    wire _556 = 1'b0;
    wire _559;
    wire _19;
    reg PHASE_5;
    wire [63:0] _640;
    wire [5:0] address_30;
    wire _590;
    wire read_enable_24;
    wire write_enable_30;
    wire _592;
    wire [5:0] address_31;
    wire _585;
    wire read_enable_25;
    wire _583;
    wire write_enable_31;
    wire _587;
    wire [131:0] _595;
    wire [63:0] _596;
    wire [63:0] _651;
    wire [63:0] data_27;
    wire [63:0] data_28;
    wire [63:0] data_29;
    wire [63:0] data_30;
    wire [5:0] address_32;
    wire _576;
    wire read_enable_26;
    wire _573;
    wire _574;
    wire write_enable_32;
    wire _578;
    wire [5:0] address_33;
    wire _569;
    wire read_enable_27;
    wire _566;
    wire _567;
    wire write_enable_33;
    wire _571;
    wire [131:0] _581;
    wire [63:0] _582;
    wire _564 = 1'b0;
    wire _563 = 1'b0;
    wire _652;
    wire _21;
    reg PHASE_6;
    wire [63:0] q0_1;
    wire _561 = 1'b0;
    wire _560 = 1'b0;
    reg _562;
    wire [63:0] _641;
    wire [191:0] _650;
    wire [63:0] _653;
    wire [63:0] data_31;
    wire [63:0] data_32;
    wire [63:0] data_33;
    wire [63:0] data_34;
    wire [5:0] address_34;
    wire _717;
    wire _716;
    wire read_enable_28;
    wire _710 = 1'b0;
    wire _709 = 1'b0;
    wire _707 = 1'b0;
    wire _706 = 1'b0;
    wire _704 = 1'b0;
    wire _703 = 1'b0;
    wire _701 = 1'b0;
    wire _700 = 1'b0;
    wire _698 = 1'b0;
    wire _697 = 1'b0;
    wire _695 = 1'b0;
    wire _694 = 1'b0;
    wire _692 = 1'b0;
    wire _691 = 1'b0;
    wire _689 = 1'b0;
    wire _688 = 1'b0;
    wire _686 = 1'b0;
    wire _685 = 1'b0;
    reg _687;
    reg _690;
    reg _693;
    reg _696;
    reg _699;
    reg _702;
    reg _705;
    reg _708;
    reg _711;
    wire _712;
    wire _683 = 1'b0;
    wire _682 = 1'b0;
    wire _680 = 1'b0;
    wire _679 = 1'b0;
    wire _677 = 1'b0;
    wire _676 = 1'b0;
    wire _674 = 1'b0;
    wire _673 = 1'b0;
    wire _671 = 1'b0;
    wire _670 = 1'b0;
    wire _668 = 1'b0;
    wire _667 = 1'b0;
    wire _665 = 1'b0;
    wire _664 = 1'b0;
    wire _662 = 1'b0;
    wire _661 = 1'b0;
    wire _659 = 1'b0;
    wire _658 = 1'b0;
    reg _660;
    reg _663;
    reg _666;
    reg _669;
    reg _672;
    reg _675;
    reg _678;
    reg _681;
    reg _684;
    wire _713;
    wire _714;
    wire write_enable_34;
    wire _719;
    wire [131:0] _726;
    wire [63:0] _727;
    wire _655 = 1'b0;
    wire _654 = 1'b0;
    wire _657;
    wire _23;
    reg PHASE_7;
    wire [63:0] _739;
    wire [5:0] address_35;
    wire write_enable_35;
    wire [5:0] address_36;
    wire _914;
    wire read_enable_29;
    wire _912;
    wire write_enable_36;
    wire _916;
    wire [131:0] _921;
    wire [63:0] _922;
    wire [5:0] _907 = 6'b000000;
    wire [5:0] address_37;
    wire _905;
    wire write_enable_37;
    wire [63:0] _830;
    wire [63:0] _829;
    wire [63:0] _831;
    wire [63:0] _827;
    wire [63:0] _826;
    wire [63:0] q1_2;
    wire [63:0] _832;
    wire [5:0] address_38;
    wire write_enable_38 = 1'b0;
    wire _817;
    wire read_enable_30;
    wire [5:0] address_39;
    wire _813;
    wire read_enable_31;
    wire _811;
    wire write_enable_39;
    wire _815;
    wire [131:0] _822;
    wire [63:0] _823;
    wire [63:0] data_35 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_36;
    wire [5:0] _805 = 6'b000000;
    wire _803;
    wire _802;
    wire _801;
    wire _800;
    wire _799;
    wire _798;
    wire [5:0] _804;
    wire [5:0] address_40;
    wire write_enable_40 = 1'b0;
    wire _795;
    wire read_enable_32;
    wire [63:0] data_37;
    wire [63:0] data_38;
    wire _792;
    wire _791;
    wire _790;
    wire _789;
    wire _788;
    wire _787;
    wire [5:0] _793;
    wire [5:0] address_41;
    wire _784;
    wire read_enable_33;
    wire _782;
    wire write_enable_41;
    wire _786;
    wire [131:0] _809;
    wire [63:0] _810;
    wire _741 = 1'b0;
    wire _740 = 1'b0;
    wire _743;
    wire _27;
    reg PHASE_8;
    wire [63:0] _824;
    wire [5:0] address_42;
    wire _774;
    wire read_enable_34;
    wire write_enable_42;
    wire _776;
    wire [5:0] address_43;
    wire _769;
    wire read_enable_35;
    wire _767;
    wire write_enable_43;
    wire _771;
    wire [131:0] _779;
    wire [63:0] _780;
    wire [63:0] _835;
    wire [63:0] data_39;
    wire [63:0] data_40;
    wire [63:0] data_41;
    wire [63:0] data_42;
    wire [5:0] address_44;
    wire _760;
    wire read_enable_36;
    wire _757;
    wire _758;
    wire write_enable_44;
    wire _762;
    wire [5:0] address_45;
    wire _753;
    wire read_enable_37;
    wire _750;
    wire _751;
    wire write_enable_45;
    wire _755;
    wire [131:0] _765;
    wire [63:0] _766;
    wire _748 = 1'b0;
    wire _747 = 1'b0;
    wire _836;
    wire _29;
    reg PHASE_9;
    wire [63:0] q0_2;
    wire _745 = 1'b0;
    wire _744 = 1'b0;
    reg _746;
    wire [63:0] _825;
    wire [191:0] _834;
    wire [63:0] _837;
    wire [63:0] data_43;
    wire [63:0] data_44;
    wire [63:0] data_45;
    wire [63:0] data_46;
    wire [5:0] address_46;
    wire _901;
    wire _900;
    wire read_enable_38;
    wire _894 = 1'b0;
    wire _893 = 1'b0;
    wire _891 = 1'b0;
    wire _890 = 1'b0;
    wire _888 = 1'b0;
    wire _887 = 1'b0;
    wire _885 = 1'b0;
    wire _884 = 1'b0;
    wire _882 = 1'b0;
    wire _881 = 1'b0;
    wire _879 = 1'b0;
    wire _878 = 1'b0;
    wire _876 = 1'b0;
    wire _875 = 1'b0;
    wire _873 = 1'b0;
    wire _872 = 1'b0;
    wire _870 = 1'b0;
    wire _869 = 1'b0;
    reg _871;
    reg _874;
    reg _877;
    reg _880;
    reg _883;
    reg _886;
    reg _889;
    reg _892;
    reg _895;
    wire _896;
    wire _867 = 1'b0;
    wire _866 = 1'b0;
    wire _864 = 1'b0;
    wire _863 = 1'b0;
    wire _861 = 1'b0;
    wire _860 = 1'b0;
    wire _858 = 1'b0;
    wire _857 = 1'b0;
    wire _855 = 1'b0;
    wire _854 = 1'b0;
    wire _852 = 1'b0;
    wire _851 = 1'b0;
    wire _849 = 1'b0;
    wire _848 = 1'b0;
    wire _846 = 1'b0;
    wire _845 = 1'b0;
    wire _843 = 1'b0;
    wire _842 = 1'b0;
    reg _844;
    reg _847;
    reg _850;
    reg _853;
    reg _856;
    reg _859;
    reg _862;
    reg _865;
    reg _868;
    wire _897;
    wire _898;
    wire write_enable_46;
    wire _903;
    wire [131:0] _910;
    wire [63:0] _911;
    wire _839 = 1'b0;
    wire _838 = 1'b0;
    wire _841;
    wire _31;
    reg PHASE_10;
    wire [63:0] _923;
    wire [5:0] address_47;
    wire write_enable_47;
    wire [5:0] address_48;
    wire _1098;
    wire read_enable_39;
    wire _1096;
    wire write_enable_48;
    wire _1100;
    wire [131:0] _1105;
    wire [63:0] _1106;
    wire [5:0] _1091 = 6'b000000;
    wire [5:0] address_49;
    wire _1089;
    wire write_enable_49;
    wire [63:0] _1014;
    wire [63:0] _1013;
    wire [63:0] _1015;
    wire [63:0] _1011;
    wire [63:0] _1010;
    wire [63:0] q1_3;
    wire [63:0] _1016;
    wire [5:0] address_50;
    wire write_enable_50 = 1'b0;
    wire _1001;
    wire read_enable_40;
    wire [5:0] address_51;
    wire _997;
    wire read_enable_41;
    wire _995;
    wire write_enable_51;
    wire _999;
    wire [131:0] _1006;
    wire [63:0] _1007;
    wire [63:0] data_47 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_48;
    wire [5:0] _989 = 6'b000000;
    wire _987;
    wire _986;
    wire _985;
    wire _984;
    wire _983;
    wire _982;
    wire [5:0] _988;
    wire [5:0] address_52;
    wire write_enable_52 = 1'b0;
    wire _979;
    wire read_enable_42;
    wire [63:0] data_49;
    wire [63:0] data_50;
    wire _976;
    wire _975;
    wire _974;
    wire _973;
    wire _972;
    wire _971;
    wire [5:0] _977;
    wire [5:0] address_53;
    wire _968;
    wire read_enable_43;
    wire _966;
    wire write_enable_53;
    wire _970;
    wire [131:0] _993;
    wire [63:0] _994;
    wire _925 = 1'b0;
    wire _924 = 1'b0;
    wire _927;
    wire _35;
    reg PHASE_11;
    wire [63:0] _1008;
    wire [5:0] address_54;
    wire _958;
    wire read_enable_44;
    wire write_enable_54;
    wire _960;
    wire [5:0] address_55;
    wire _953;
    wire read_enable_45;
    wire _951;
    wire write_enable_55;
    wire _955;
    wire [131:0] _963;
    wire [63:0] _964;
    wire [63:0] _1019;
    wire [63:0] data_51;
    wire [63:0] data_52;
    wire [63:0] data_53;
    wire [63:0] data_54;
    wire [5:0] address_56;
    wire _944;
    wire read_enable_46;
    wire _941;
    wire _942;
    wire write_enable_56;
    wire _946;
    wire [5:0] address_57;
    wire _937;
    wire read_enable_47;
    wire _934;
    wire _935;
    wire write_enable_57;
    wire _939;
    wire [131:0] _949;
    wire [63:0] _950;
    wire _932 = 1'b0;
    wire _931 = 1'b0;
    wire _1020;
    wire _37;
    reg PHASE_12;
    wire [63:0] q0_3;
    wire _929 = 1'b0;
    wire _928 = 1'b0;
    reg _930;
    wire [63:0] _1009;
    wire [191:0] _1018;
    wire [63:0] _1021;
    wire [63:0] data_55;
    wire [63:0] data_56;
    wire [63:0] data_57;
    wire [63:0] data_58;
    wire [5:0] address_58;
    wire _1085;
    wire _1084;
    wire read_enable_48;
    wire _1078 = 1'b0;
    wire _1077 = 1'b0;
    wire _1075 = 1'b0;
    wire _1074 = 1'b0;
    wire _1072 = 1'b0;
    wire _1071 = 1'b0;
    wire _1069 = 1'b0;
    wire _1068 = 1'b0;
    wire _1066 = 1'b0;
    wire _1065 = 1'b0;
    wire _1063 = 1'b0;
    wire _1062 = 1'b0;
    wire _1060 = 1'b0;
    wire _1059 = 1'b0;
    wire _1057 = 1'b0;
    wire _1056 = 1'b0;
    wire _1054 = 1'b0;
    wire _1053 = 1'b0;
    reg _1055;
    reg _1058;
    reg _1061;
    reg _1064;
    reg _1067;
    reg _1070;
    reg _1073;
    reg _1076;
    reg _1079;
    wire _1080;
    wire _1051 = 1'b0;
    wire _1050 = 1'b0;
    wire _1048 = 1'b0;
    wire _1047 = 1'b0;
    wire _1045 = 1'b0;
    wire _1044 = 1'b0;
    wire _1042 = 1'b0;
    wire _1041 = 1'b0;
    wire _1039 = 1'b0;
    wire _1038 = 1'b0;
    wire _1036 = 1'b0;
    wire _1035 = 1'b0;
    wire _1033 = 1'b0;
    wire _1032 = 1'b0;
    wire _1030 = 1'b0;
    wire _1029 = 1'b0;
    wire _1027 = 1'b0;
    wire _1026 = 1'b0;
    reg _1028;
    reg _1031;
    reg _1034;
    reg _1037;
    reg _1040;
    reg _1043;
    reg _1046;
    reg _1049;
    reg _1052;
    wire _1081;
    wire _1082;
    wire write_enable_58;
    wire _1087;
    wire [131:0] _1094;
    wire [63:0] _1095;
    wire _1023 = 1'b0;
    wire _1022 = 1'b0;
    wire _1025;
    wire _39;
    reg PHASE_13;
    wire [63:0] _1107;
    wire [5:0] address_59;
    wire write_enable_59;
    wire [5:0] address_60;
    wire _1282;
    wire read_enable_49;
    wire _1280;
    wire write_enable_60;
    wire _1284;
    wire [131:0] _1289;
    wire [63:0] _1290;
    wire [5:0] _1275 = 6'b000000;
    wire [5:0] address_61;
    wire _1273;
    wire write_enable_61;
    wire [63:0] _1198;
    wire [63:0] _1197;
    wire [63:0] _1199;
    wire [63:0] _1195;
    wire [63:0] _1194;
    wire [63:0] q1_4;
    wire [63:0] _1200;
    wire [5:0] address_62;
    wire write_enable_62 = 1'b0;
    wire _1185;
    wire read_enable_50;
    wire [5:0] address_63;
    wire _1181;
    wire read_enable_51;
    wire _1179;
    wire write_enable_63;
    wire _1183;
    wire [131:0] _1190;
    wire [63:0] _1191;
    wire [63:0] data_59 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_60;
    wire [5:0] _1173 = 6'b000000;
    wire _1171;
    wire _1170;
    wire _1169;
    wire _1168;
    wire _1167;
    wire _1166;
    wire [5:0] _1172;
    wire [5:0] address_64;
    wire write_enable_64 = 1'b0;
    wire _1163;
    wire read_enable_52;
    wire [63:0] data_61;
    wire [63:0] data_62;
    wire _1160;
    wire _1159;
    wire _1158;
    wire _1157;
    wire _1156;
    wire _1155;
    wire [5:0] _1161;
    wire [5:0] address_65;
    wire _1152;
    wire read_enable_53;
    wire _1150;
    wire write_enable_65;
    wire _1154;
    wire [131:0] _1177;
    wire [63:0] _1178;
    wire _1109 = 1'b0;
    wire _1108 = 1'b0;
    wire _1111;
    wire _43;
    reg PHASE_14;
    wire [63:0] _1192;
    wire [5:0] address_66;
    wire _1142;
    wire read_enable_54;
    wire write_enable_66;
    wire _1144;
    wire [5:0] address_67;
    wire _1137;
    wire read_enable_55;
    wire _1135;
    wire write_enable_67;
    wire _1139;
    wire [131:0] _1147;
    wire [63:0] _1148;
    wire [63:0] _1203;
    wire [63:0] data_63;
    wire [63:0] data_64;
    wire [63:0] data_65;
    wire [63:0] data_66;
    wire [5:0] address_68;
    wire _1128;
    wire read_enable_56;
    wire _1125;
    wire _1126;
    wire write_enable_68;
    wire _1130;
    wire [5:0] address_69;
    wire _1121;
    wire read_enable_57;
    wire _1118;
    wire _1119;
    wire write_enable_69;
    wire _1123;
    wire [131:0] _1133;
    wire [63:0] _1134;
    wire _1116 = 1'b0;
    wire _1115 = 1'b0;
    wire _1204;
    wire _45;
    reg PHASE_15;
    wire [63:0] q0_4;
    wire _1113 = 1'b0;
    wire _1112 = 1'b0;
    reg _1114;
    wire [63:0] _1193;
    wire [191:0] _1202;
    wire [63:0] _1205;
    wire [63:0] data_67;
    wire [63:0] data_68;
    wire [63:0] data_69;
    wire [63:0] data_70;
    wire [5:0] address_70;
    wire _1269;
    wire _1268;
    wire read_enable_58;
    wire _1262 = 1'b0;
    wire _1261 = 1'b0;
    wire _1259 = 1'b0;
    wire _1258 = 1'b0;
    wire _1256 = 1'b0;
    wire _1255 = 1'b0;
    wire _1253 = 1'b0;
    wire _1252 = 1'b0;
    wire _1250 = 1'b0;
    wire _1249 = 1'b0;
    wire _1247 = 1'b0;
    wire _1246 = 1'b0;
    wire _1244 = 1'b0;
    wire _1243 = 1'b0;
    wire _1241 = 1'b0;
    wire _1240 = 1'b0;
    wire _1238 = 1'b0;
    wire _1237 = 1'b0;
    reg _1239;
    reg _1242;
    reg _1245;
    reg _1248;
    reg _1251;
    reg _1254;
    reg _1257;
    reg _1260;
    reg _1263;
    wire _1264;
    wire _1235 = 1'b0;
    wire _1234 = 1'b0;
    wire _1232 = 1'b0;
    wire _1231 = 1'b0;
    wire _1229 = 1'b0;
    wire _1228 = 1'b0;
    wire _1226 = 1'b0;
    wire _1225 = 1'b0;
    wire _1223 = 1'b0;
    wire _1222 = 1'b0;
    wire _1220 = 1'b0;
    wire _1219 = 1'b0;
    wire _1217 = 1'b0;
    wire _1216 = 1'b0;
    wire _1214 = 1'b0;
    wire _1213 = 1'b0;
    wire _1211 = 1'b0;
    wire _1210 = 1'b0;
    reg _1212;
    reg _1215;
    reg _1218;
    reg _1221;
    reg _1224;
    reg _1227;
    reg _1230;
    reg _1233;
    reg _1236;
    wire _1265;
    wire _1266;
    wire write_enable_70;
    wire _1271;
    wire [131:0] _1278;
    wire [63:0] _1279;
    wire _1207 = 1'b0;
    wire _1206 = 1'b0;
    wire _1209;
    wire _47;
    reg PHASE_16;
    wire [63:0] _1291;
    wire [5:0] address_71;
    wire write_enable_71;
    wire [5:0] address_72;
    wire _1466;
    wire read_enable_59;
    wire _1464;
    wire write_enable_72;
    wire _1468;
    wire [131:0] _1473;
    wire [63:0] _1474;
    wire [5:0] _1459 = 6'b000000;
    wire [5:0] address_73;
    wire _1457;
    wire write_enable_73;
    wire [63:0] _1382;
    wire [63:0] _1381;
    wire [63:0] _1383;
    wire [63:0] _1379;
    wire [63:0] _1378;
    wire [63:0] q1_5;
    wire [63:0] _1384;
    wire [5:0] address_74;
    wire write_enable_74 = 1'b0;
    wire _1369;
    wire read_enable_60;
    wire [5:0] address_75;
    wire _1365;
    wire read_enable_61;
    wire _1363;
    wire write_enable_75;
    wire _1367;
    wire [131:0] _1374;
    wire [63:0] _1375;
    wire [63:0] data_71 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_72;
    wire [5:0] _1357 = 6'b000000;
    wire _1355;
    wire _1354;
    wire _1353;
    wire _1352;
    wire _1351;
    wire _1350;
    wire [5:0] _1356;
    wire [5:0] address_76;
    wire write_enable_76 = 1'b0;
    wire _1347;
    wire read_enable_62;
    wire [63:0] data_73;
    wire [63:0] data_74;
    wire _1344;
    wire _1343;
    wire _1342;
    wire _1341;
    wire _1340;
    wire _1339;
    wire [5:0] _1345;
    wire [5:0] address_77;
    wire _1336;
    wire read_enable_63;
    wire _1334;
    wire write_enable_77;
    wire _1338;
    wire [131:0] _1361;
    wire [63:0] _1362;
    wire _1293 = 1'b0;
    wire _1292 = 1'b0;
    wire _1295;
    wire _51;
    reg PHASE_17;
    wire [63:0] _1376;
    wire [5:0] address_78;
    wire _1326;
    wire read_enable_64;
    wire write_enable_78;
    wire _1328;
    wire [5:0] address_79;
    wire _1321;
    wire read_enable_65;
    wire _1319;
    wire write_enable_79;
    wire _1323;
    wire [131:0] _1331;
    wire [63:0] _1332;
    wire [63:0] _1387;
    wire [63:0] data_75;
    wire [63:0] data_76;
    wire [63:0] data_77;
    wire [63:0] data_78;
    wire [5:0] address_80;
    wire _1312;
    wire read_enable_66;
    wire _1309;
    wire _1310;
    wire write_enable_80;
    wire _1314;
    wire [5:0] address_81;
    wire _1305;
    wire read_enable_67;
    wire _1302;
    wire _1303;
    wire write_enable_81;
    wire _1307;
    wire [131:0] _1317;
    wire [63:0] _1318;
    wire _1300 = 1'b0;
    wire _1299 = 1'b0;
    wire _1388;
    wire _53;
    reg PHASE_18;
    wire [63:0] q0_5;
    wire _1297 = 1'b0;
    wire _1296 = 1'b0;
    reg _1298;
    wire [63:0] _1377;
    wire [191:0] _1386;
    wire [63:0] _1389;
    wire [63:0] data_79;
    wire [63:0] data_80;
    wire [63:0] data_81;
    wire [63:0] data_82;
    wire [5:0] address_82;
    wire _1453;
    wire _1452;
    wire read_enable_68;
    wire _1446 = 1'b0;
    wire _1445 = 1'b0;
    wire _1443 = 1'b0;
    wire _1442 = 1'b0;
    wire _1440 = 1'b0;
    wire _1439 = 1'b0;
    wire _1437 = 1'b0;
    wire _1436 = 1'b0;
    wire _1434 = 1'b0;
    wire _1433 = 1'b0;
    wire _1431 = 1'b0;
    wire _1430 = 1'b0;
    wire _1428 = 1'b0;
    wire _1427 = 1'b0;
    wire _1425 = 1'b0;
    wire _1424 = 1'b0;
    wire _1422 = 1'b0;
    wire _1421 = 1'b0;
    reg _1423;
    reg _1426;
    reg _1429;
    reg _1432;
    reg _1435;
    reg _1438;
    reg _1441;
    reg _1444;
    reg _1447;
    wire _1448;
    wire _1419 = 1'b0;
    wire _1418 = 1'b0;
    wire _1416 = 1'b0;
    wire _1415 = 1'b0;
    wire _1413 = 1'b0;
    wire _1412 = 1'b0;
    wire _1410 = 1'b0;
    wire _1409 = 1'b0;
    wire _1407 = 1'b0;
    wire _1406 = 1'b0;
    wire _1404 = 1'b0;
    wire _1403 = 1'b0;
    wire _1401 = 1'b0;
    wire _1400 = 1'b0;
    wire _1398 = 1'b0;
    wire _1397 = 1'b0;
    wire _1395 = 1'b0;
    wire _1394 = 1'b0;
    reg _1396;
    reg _1399;
    reg _1402;
    reg _1405;
    reg _1408;
    reg _1411;
    reg _1414;
    reg _1417;
    reg _1420;
    wire _1449;
    wire _1450;
    wire write_enable_82;
    wire _1455;
    wire [131:0] _1462;
    wire [63:0] _1463;
    wire _1391 = 1'b0;
    wire _1390 = 1'b0;
    wire _1393;
    wire _55;
    reg PHASE_19;
    wire [63:0] _1475;
    wire [5:0] address_83;
    wire write_enable_83;
    wire [5:0] address_84;
    wire _1650;
    wire read_enable_69;
    wire _1648;
    wire write_enable_84;
    wire _1652;
    wire [131:0] _1657;
    wire [63:0] _1658;
    wire [5:0] _1643 = 6'b000000;
    wire [5:0] address_85;
    wire _1641;
    wire write_enable_85;
    wire [3:0] _280;
    wire _279;
    wire _277;
    wire [63:0] _276;
    wire [63:0] _275;
    wire [63:0] _274;
    wire [63:0] _273;
    wire [63:0] _272;
    wire [63:0] _271;
    wire [63:0] _270;
    wire [63:0] _1566;
    wire [63:0] _1565;
    wire [63:0] _1567;
    wire [63:0] _1563;
    wire [63:0] _1562;
    wire [63:0] q1_6;
    wire [63:0] _1568;
    wire [5:0] address_86;
    wire write_enable_86 = 1'b0;
    wire _1553;
    wire read_enable_70;
    wire [5:0] address_87;
    wire _1549;
    wire read_enable_71;
    wire _1547;
    wire write_enable_87;
    wire _1551;
    wire [131:0] _1558;
    wire [63:0] _1559;
    wire [63:0] data_83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_84;
    wire [5:0] _1541 = 6'b000000;
    wire _1539;
    wire _1538;
    wire _1537;
    wire _1536;
    wire _1535;
    wire _1534;
    wire [5:0] _1540;
    wire [5:0] address_88;
    wire write_enable_88 = 1'b0;
    wire _1531;
    wire read_enable_72;
    wire [63:0] data_85;
    wire [63:0] data_86;
    wire [5:0] _60;
    wire _1528;
    wire _1527;
    wire _1526;
    wire _1525;
    wire _1524;
    wire _1523;
    wire [5:0] _1529;
    wire [5:0] address_89;
    wire _1520;
    wire read_enable_73;
    wire [7:0] _62;
    wire _1518;
    wire write_enable_89;
    wire _1522;
    wire [131:0] _1545;
    wire [63:0] _1546;
    wire _1477 = 1'b0;
    wire _1476 = 1'b0;
    wire _1479;
    wire _63;
    reg PHASE_20;
    wire [63:0] _1560;
    wire [5:0] address_90;
    wire _1510;
    wire read_enable_74;
    wire write_enable_90;
    wire _1512;
    wire [5:0] address_91;
    wire _1505;
    wire read_enable_75;
    wire _1503;
    wire write_enable_91;
    wire _1507;
    wire [131:0] _1515;
    wire [63:0] _1516;
    wire [63:0] _1571;
    wire [63:0] data_87;
    wire [63:0] data_88;
    wire [63:0] data_89;
    wire [63:0] data_90;
    wire [5:0] _198 = 6'b000000;
    wire [5:0] _197 = 6'b000000;
    wire [5:0] _195 = 6'b000000;
    wire [5:0] _194 = 6'b000000;
    wire [5:0] _192 = 6'b000000;
    wire [5:0] _191 = 6'b000000;
    wire [5:0] _189 = 6'b000000;
    wire [5:0] _188 = 6'b000000;
    wire [5:0] _186 = 6'b000000;
    wire [5:0] _185 = 6'b000000;
    wire [5:0] _183 = 6'b000000;
    wire [5:0] _182 = 6'b000000;
    wire [5:0] _180 = 6'b000000;
    wire [5:0] _179 = 6'b000000;
    wire [5:0] _177 = 6'b000000;
    wire [5:0] _176 = 6'b000000;
    wire [5:0] _174 = 6'b000000;
    wire [5:0] _173 = 6'b000000;
    reg [5:0] _175;
    reg [5:0] _178;
    reg [5:0] _181;
    reg [5:0] _184;
    reg [5:0] _187;
    reg [5:0] _190;
    reg [5:0] _193;
    reg [5:0] _196;
    reg [5:0] _199;
    wire [5:0] _172;
    wire [5:0] address_92;
    wire _1496;
    wire read_enable_76;
    wire _1493;
    wire _1494;
    wire write_enable_92;
    wire _1498;
    wire [5:0] address_93;
    wire _1489;
    wire read_enable_77;
    wire _1486;
    wire _1487;
    wire write_enable_93;
    wire _1491;
    wire [131:0] _1501;
    wire [63:0] _1502;
    wire _99;
    wire _1484 = 1'b0;
    wire _1483 = 1'b0;
    wire _1572;
    wire _65;
    reg PHASE_21;
    wire [63:0] q0_6;
    wire _1481 = 1'b0;
    wire _1480 = 1'b0;
    wire _92;
    reg _1482;
    wire [63:0] _1561;
    wire [191:0] _1570;
    wire [63:0] _1573;
    wire [63:0] data_91;
    wire [63:0] data_92;
    wire [63:0] data_93;
    wire [63:0] data_94;
    wire [5:0] _163 = 6'b000000;
    wire [5:0] _162 = 6'b000000;
    wire [5:0] _160 = 6'b000000;
    wire [5:0] _159 = 6'b000000;
    wire [5:0] _157 = 6'b000000;
    wire [5:0] _156 = 6'b000000;
    wire [5:0] _154 = 6'b000000;
    wire [5:0] _153 = 6'b000000;
    wire [5:0] _151 = 6'b000000;
    wire [5:0] _150 = 6'b000000;
    wire [5:0] _148 = 6'b000000;
    wire [5:0] _147 = 6'b000000;
    wire [5:0] _145 = 6'b000000;
    wire [5:0] _144 = 6'b000000;
    wire [5:0] _142 = 6'b000000;
    wire [5:0] _141 = 6'b000000;
    wire [5:0] _139 = 6'b000000;
    wire [5:0] _138 = 6'b000000;
    wire [5:0] _137;
    reg [5:0] _140;
    reg [5:0] _143;
    reg [5:0] _146;
    reg [5:0] _149;
    reg [5:0] _152;
    reg [5:0] _155;
    reg [5:0] _158;
    reg [5:0] _161;
    reg [5:0] _164;
    wire [5:0] _68;
    wire [5:0] address_94;
    wire _1637;
    wire [7:0] _70;
    wire _1636;
    wire read_enable_78;
    wire _1630 = 1'b0;
    wire _1629 = 1'b0;
    wire _1627 = 1'b0;
    wire _1626 = 1'b0;
    wire _1624 = 1'b0;
    wire _1623 = 1'b0;
    wire _1621 = 1'b0;
    wire _1620 = 1'b0;
    wire _1618 = 1'b0;
    wire _1617 = 1'b0;
    wire _1615 = 1'b0;
    wire _1614 = 1'b0;
    wire _1612 = 1'b0;
    wire _1611 = 1'b0;
    wire _1609 = 1'b0;
    wire _1608 = 1'b0;
    wire _1606 = 1'b0;
    wire _1605 = 1'b0;
    wire _278;
    reg _1607;
    reg _1610;
    reg _1613;
    reg _1616;
    reg _1619;
    reg _1622;
    reg _1625;
    reg _1628;
    reg _1631;
    wire _1632;
    wire _1603 = 1'b0;
    wire _1602 = 1'b0;
    wire _1600 = 1'b0;
    wire _1599 = 1'b0;
    wire _1597 = 1'b0;
    wire _1596 = 1'b0;
    wire _1594 = 1'b0;
    wire _1593 = 1'b0;
    wire _1591 = 1'b0;
    wire _1590 = 1'b0;
    wire _1588 = 1'b0;
    wire _1587 = 1'b0;
    wire _1585 = 1'b0;
    wire _1584 = 1'b0;
    wire _1582 = 1'b0;
    wire _1581 = 1'b0;
    wire _1579 = 1'b0;
    wire _1578 = 1'b0;
    wire _130;
    reg _1580;
    reg _1583;
    reg _1586;
    reg _1589;
    reg _1592;
    reg _1595;
    reg _1598;
    reg _1601;
    reg _1604;
    wire _1633;
    wire _128 = 1'b0;
    wire _127 = 1'b0;
    wire _125 = 1'b0;
    wire _124 = 1'b0;
    wire _122 = 1'b0;
    wire _121 = 1'b0;
    wire _119 = 1'b0;
    wire _118 = 1'b0;
    wire _116 = 1'b0;
    wire _115 = 1'b0;
    wire _113 = 1'b0;
    wire _112 = 1'b0;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire vdd = 1'b1;
    wire _104 = 1'b0;
    wire _103 = 1'b0;
    wire _102;
    reg _105;
    reg _108;
    reg _111;
    reg _114;
    reg _117;
    reg _120;
    reg _123;
    reg _126;
    reg _129;
    wire _1634;
    wire write_enable_94;
    wire _1639;
    wire gnd = 1'b0;
    wire [131:0] _1646;
    wire [63:0] _1647;
    wire _72;
    wire _1575 = 1'b0;
    wire _1574 = 1'b0;
    wire _1577;
    wire _73;
    reg PHASE_22;
    wire [63:0] _1659;
    wire _76;
    wire _78;
    wire _80;
    wire _82;
    wire _84;
    wire [492:0] _91;
    wire _1660;

    /* logic */
    assign address = _360 ? _199 : _355;
    assign write_enable = _353 & _360;
    assign address_0 = _360 ? _164 : _68;
    assign _362 = ~ _360;
    assign read_enable = _348 & _362;
    assign _360 = ~ PHASE_1;
    assign write_enable_0 = _346 & _360;
    assign _364 = write_enable_0 | read_enable;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_364), .regcea(vdd), .wea(write_enable_0), .addra(address_0), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable), .regceb(vdd), .web(write_enable), .addrb(address), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_369[131:131]), .sbiterrb(_369[130:130]), .doutb(_369[129:66]), .dbiterra(_369[65:65]), .sbiterra(_369[64:64]), .douta(_369[63:0]) );
    assign _370 = _369[63:0];
    assign address_1 = PHASE_1 ? _199 : _355;
    assign _353 = _129 & _316;
    assign write_enable_1 = _353 & PHASE_1;
    assign _267 = _259[129:66];
    assign _266 = _246[129:66];
    assign _268 = PHASE ? _267 : _266;
    assign _264 = _216[129:66];
    assign _263 = _202[129:66];
    assign q1 = PHASE_0 ? _264 : _263;
    assign _269 = _96 ? _268 : q1;
    assign address_2 = _248 ? _242 : _241;
    assign _254 = ~ _248;
    assign read_enable_0 = _102 & _254;
    assign address_3 = _248 ? _60 : _230;
    assign _250 = ~ _248;
    assign read_enable_1 = _102 & _250;
    assign _248 = ~ PHASE;
    assign write_enable_3 = _219 & _248;
    assign _252 = write_enable_3 | read_enable_1;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_0
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_252), .regcea(vdd), .wea(write_enable_3), .addra(address_3), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_0), .regceb(vdd), .web(write_enable_2), .addrb(address_2), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_259[131:131]), .sbiterrb(_259[130:130]), .doutb(_259[129:66]), .dbiterra(_259[65:65]), .sbiterra(_259[64:64]), .douta(_259[63:0]) );
    assign _260 = _259[63:0];
    assign _240 = _172[5:5];
    assign _239 = _172[4:4];
    assign _238 = _172[3:3];
    assign _237 = _172[2:2];
    assign _236 = _172[1:1];
    assign _235 = _172[0:0];
    assign _241 = { _235, _236, _237, _238, _239, _240 };
    assign address_4 = PHASE ? _242 : _241;
    assign _232 = ~ PHASE;
    assign read_enable_2 = _102 & _232;
    assign data_1 = wr_d7;
    assign _229 = _137[5:5];
    assign _228 = _137[4:4];
    assign _227 = _137[3:3];
    assign _226 = _137[2:2];
    assign _225 = _137[1:1];
    assign _224 = _137[0:0];
    assign _230 = { _224, _225, _226, _227, _228, _229 };
    assign address_5 = PHASE ? _60 : _230;
    assign _221 = ~ PHASE;
    assign read_enable_3 = _102 & _221;
    assign _219 = _62[7:7];
    assign write_enable_5 = _219 & PHASE;
    assign _223 = write_enable_5 | read_enable_3;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_1
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_223), .regcea(vdd), .wea(write_enable_5), .addra(address_5), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_2), .regceb(vdd), .web(write_enable_4), .addrb(address_4), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_246[131:131]), .sbiterrb(_246[130:130]), .doutb(_246[129:66]), .dbiterra(_246[65:65]), .sbiterra(_246[64:64]), .douta(_246[63:0]) );
    assign _247 = _246[63:0];
    assign _89 = ~ PHASE;
    assign _3 = _89;
    always @(posedge _84) begin
        if (_82)
            PHASE <= _87;
        else
            if (_72)
                PHASE <= _3;
    end
    assign _261 = PHASE ? _260 : _247;
    assign address_6 = _204 ? _199 : _172;
    assign _211 = ~ _204;
    assign read_enable_4 = _102 & _211;
    assign write_enable_6 = _167 & _204;
    assign _213 = write_enable_6 | read_enable_4;
    assign address_7 = _204 ? _164 : _137;
    assign _206 = ~ _204;
    assign read_enable_5 = _102 & _206;
    assign _204 = ~ PHASE_0;
    assign write_enable_7 = _132 & _204;
    assign _208 = write_enable_7 | read_enable_5;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_2
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_208), .regcea(vdd), .wea(write_enable_7), .addra(address_7), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_213), .regceb(vdd), .web(write_enable_6), .addrb(address_6), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_216[131:131]), .sbiterrb(_216[130:130]), .doutb(_216[129:66]), .dbiterra(_216[65:65]), .sbiterra(_216[64:64]), .douta(_216[63:0]) );
    assign _217 = _216[63:0];
    assign _283 = _282[127:64];
    assign data_3 = _283;
    assign address_8 = PHASE_0 ? _199 : _172;
    assign _169 = ~ PHASE_0;
    assign read_enable_6 = _102 & _169;
    assign _166 = ~ _130;
    assign _167 = _129 & _166;
    assign write_enable_8 = _167 & PHASE_0;
    assign _171 = write_enable_8 | read_enable_6;
    assign address_9 = PHASE_0 ? _164 : _137;
    assign _134 = ~ PHASE_0;
    assign read_enable_7 = _102 & _134;
    assign _131 = ~ _130;
    assign _132 = _129 & _131;
    assign write_enable_9 = _132 & PHASE_0;
    assign _136 = write_enable_9 | read_enable_7;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_3
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_136), .regcea(vdd), .wea(write_enable_9), .addra(address_9), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_171), .regceb(vdd), .web(write_enable_8), .addrb(address_8), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_202[131:131]), .sbiterrb(_202[130:130]), .doutb(_202[129:66]), .dbiterra(_202[65:65]), .sbiterra(_202[64:64]), .douta(_202[63:0]) );
    assign _203 = _202[63:0];
    assign _284 = ~ PHASE_0;
    assign _5 = _284;
    always @(posedge _84) begin
        if (_82)
            PHASE_0 <= _98;
        else
            if (_99)
                PHASE_0 <= _5;
    end
    assign q0 = PHASE_0 ? _217 : _203;
    always @(posedge _84) begin
        if (_82)
            _96 <= _94;
        else
            _96 <= _92;
    end
    assign _262 = _96 ? _261 : q0;
    dp_14
        dp_6
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_262), .d2(_269), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_282[191:128]), .q2(_282[127:64]), .q1(_282[63:0]) );
    assign _285 = _282[63:0];
    assign data_7 = _285;
    assign address_10 = PHASE_1 ? _164 : _68;
    assign _349 = ~ PHASE_1;
    assign _348 = _70[7:7];
    assign read_enable_8 = _348 & _349;
    always @(posedge _84) begin
        if (_82)
            _319 <= _318;
        else
            _319 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _322 <= _321;
        else
            _322 <= _319;
    end
    always @(posedge _84) begin
        if (_82)
            _325 <= _324;
        else
            _325 <= _322;
    end
    always @(posedge _84) begin
        if (_82)
            _328 <= _327;
        else
            _328 <= _325;
    end
    always @(posedge _84) begin
        if (_82)
            _331 <= _330;
        else
            _331 <= _328;
    end
    always @(posedge _84) begin
        if (_82)
            _334 <= _333;
        else
            _334 <= _331;
    end
    always @(posedge _84) begin
        if (_82)
            _337 <= _336;
        else
            _337 <= _334;
    end
    always @(posedge _84) begin
        if (_82)
            _340 <= _339;
        else
            _340 <= _337;
    end
    always @(posedge _84) begin
        if (_82)
            _343 <= _342;
        else
            _343 <= _340;
    end
    assign _344 = ~ _343;
    always @(posedge _84) begin
        if (_82)
            _292 <= _291;
        else
            _292 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _295 <= _294;
        else
            _295 <= _292;
    end
    always @(posedge _84) begin
        if (_82)
            _298 <= _297;
        else
            _298 <= _295;
    end
    always @(posedge _84) begin
        if (_82)
            _301 <= _300;
        else
            _301 <= _298;
    end
    always @(posedge _84) begin
        if (_82)
            _304 <= _303;
        else
            _304 <= _301;
    end
    always @(posedge _84) begin
        if (_82)
            _307 <= _306;
        else
            _307 <= _304;
    end
    always @(posedge _84) begin
        if (_82)
            _310 <= _309;
        else
            _310 <= _307;
    end
    always @(posedge _84) begin
        if (_82)
            _313 <= _312;
        else
            _313 <= _310;
    end
    always @(posedge _84) begin
        if (_82)
            _316 <= _315;
        else
            _316 <= _313;
    end
    assign _345 = _316 & _344;
    assign _346 = _129 & _345;
    assign write_enable_10 = _346 & PHASE_1;
    assign _351 = write_enable_10 | read_enable_8;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_4
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_351), .regcea(vdd), .wea(write_enable_10), .addra(address_10), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_1), .regceb(vdd), .web(write_enable_1), .addrb(address_1), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_358[131:131]), .sbiterrb(_358[130:130]), .doutb(_358[129:66]), .dbiterra(_358[65:65]), .sbiterra(_358[64:64]), .douta(_358[63:0]) );
    assign _359 = _358[63:0];
    assign _289 = ~ PHASE_1;
    assign _7 = _289;
    always @(posedge _84) begin
        if (_82)
            PHASE_1 <= _287;
        else
            if (_72)
                PHASE_1 <= _7;
    end
    assign _371 = PHASE_1 ? _370 : _359;
    assign address_11 = _544 ? _199 : _539;
    assign write_enable_11 = _537 & _544;
    assign address_12 = _544 ? _164 : _68;
    assign _546 = ~ _544;
    assign read_enable_9 = _532 & _546;
    assign _544 = ~ PHASE_4;
    assign write_enable_12 = _530 & _544;
    assign _548 = write_enable_12 | read_enable_9;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_5
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_548), .regcea(vdd), .wea(write_enable_12), .addra(address_12), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_11), .regceb(vdd), .web(write_enable_11), .addrb(address_11), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_553[131:131]), .sbiterrb(_553[130:130]), .doutb(_553[129:66]), .dbiterra(_553[65:65]), .sbiterra(_553[64:64]), .douta(_553[63:0]) );
    assign _554 = _553[63:0];
    assign address_13 = PHASE_4 ? _199 : _539;
    assign _537 = _129 & _500;
    assign write_enable_13 = _537 & PHASE_4;
    assign _462 = _454[129:66];
    assign _461 = _441[129:66];
    assign _463 = PHASE_2 ? _462 : _461;
    assign _459 = _411[129:66];
    assign _458 = _397[129:66];
    assign q1_0 = PHASE_3 ? _459 : _458;
    assign _464 = _378 ? _463 : q1_0;
    assign address_14 = _443 ? _437 : _436;
    assign _449 = ~ _443;
    assign read_enable_10 = _102 & _449;
    assign address_15 = _443 ? _60 : _425;
    assign _445 = ~ _443;
    assign read_enable_11 = _102 & _445;
    assign _443 = ~ PHASE_2;
    assign write_enable_15 = _414 & _443;
    assign _447 = write_enable_15 | read_enable_11;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_6
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_447), .regcea(vdd), .wea(write_enable_15), .addra(address_15), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_10), .regceb(vdd), .web(write_enable_14), .addrb(address_14), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_454[131:131]), .sbiterrb(_454[130:130]), .doutb(_454[129:66]), .dbiterra(_454[65:65]), .sbiterra(_454[64:64]), .douta(_454[63:0]) );
    assign _455 = _454[63:0];
    assign _435 = _172[5:5];
    assign _434 = _172[4:4];
    assign _433 = _172[3:3];
    assign _432 = _172[2:2];
    assign _431 = _172[1:1];
    assign _430 = _172[0:0];
    assign _436 = { _430, _431, _432, _433, _434, _435 };
    assign address_16 = PHASE_2 ? _437 : _436;
    assign _427 = ~ PHASE_2;
    assign read_enable_12 = _102 & _427;
    assign data_13 = wr_d6;
    assign _424 = _137[5:5];
    assign _423 = _137[4:4];
    assign _422 = _137[3:3];
    assign _421 = _137[2:2];
    assign _420 = _137[1:1];
    assign _419 = _137[0:0];
    assign _425 = { _419, _420, _421, _422, _423, _424 };
    assign address_17 = PHASE_2 ? _60 : _425;
    assign _416 = ~ PHASE_2;
    assign read_enable_13 = _102 & _416;
    assign _414 = _62[6:6];
    assign write_enable_17 = _414 & PHASE_2;
    assign _418 = write_enable_17 | read_enable_13;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_7
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_418), .regcea(vdd), .wea(write_enable_17), .addra(address_17), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_12), .regceb(vdd), .web(write_enable_16), .addrb(address_16), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_441[131:131]), .sbiterrb(_441[130:130]), .doutb(_441[129:66]), .dbiterra(_441[65:65]), .sbiterra(_441[64:64]), .douta(_441[63:0]) );
    assign _442 = _441[63:0];
    assign _375 = ~ PHASE_2;
    assign _11 = _375;
    always @(posedge _84) begin
        if (_82)
            PHASE_2 <= _373;
        else
            if (_72)
                PHASE_2 <= _11;
    end
    assign _456 = PHASE_2 ? _455 : _442;
    assign address_18 = _399 ? _199 : _172;
    assign _406 = ~ _399;
    assign read_enable_14 = _102 & _406;
    assign write_enable_18 = _390 & _399;
    assign _408 = write_enable_18 | read_enable_14;
    assign address_19 = _399 ? _164 : _137;
    assign _401 = ~ _399;
    assign read_enable_15 = _102 & _401;
    assign _399 = ~ PHASE_3;
    assign write_enable_19 = _383 & _399;
    assign _403 = write_enable_19 | read_enable_15;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_8
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_403), .regcea(vdd), .wea(write_enable_19), .addra(address_19), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_408), .regceb(vdd), .web(write_enable_18), .addrb(address_18), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_411[131:131]), .sbiterrb(_411[130:130]), .doutb(_411[129:66]), .dbiterra(_411[65:65]), .sbiterra(_411[64:64]), .douta(_411[63:0]) );
    assign _412 = _411[63:0];
    assign _467 = _466[127:64];
    assign data_15 = _467;
    assign address_20 = PHASE_3 ? _199 : _172;
    assign _392 = ~ PHASE_3;
    assign read_enable_16 = _102 & _392;
    assign _389 = ~ _130;
    assign _390 = _129 & _389;
    assign write_enable_20 = _390 & PHASE_3;
    assign _394 = write_enable_20 | read_enable_16;
    assign address_21 = PHASE_3 ? _164 : _137;
    assign _385 = ~ PHASE_3;
    assign read_enable_17 = _102 & _385;
    assign _382 = ~ _130;
    assign _383 = _129 & _382;
    assign write_enable_21 = _383 & PHASE_3;
    assign _387 = write_enable_21 | read_enable_17;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_9
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_387), .regcea(vdd), .wea(write_enable_21), .addra(address_21), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_394), .regceb(vdd), .web(write_enable_20), .addrb(address_20), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_397[131:131]), .sbiterrb(_397[130:130]), .doutb(_397[129:66]), .dbiterra(_397[65:65]), .sbiterra(_397[64:64]), .douta(_397[63:0]) );
    assign _398 = _397[63:0];
    assign _468 = ~ PHASE_3;
    assign _13 = _468;
    always @(posedge _84) begin
        if (_82)
            PHASE_3 <= _380;
        else
            if (_99)
                PHASE_3 <= _13;
    end
    assign q0_0 = PHASE_3 ? _412 : _398;
    always @(posedge _84) begin
        if (_82)
            _378 <= _377;
        else
            _378 <= _92;
    end
    assign _457 = _378 ? _456 : q0_0;
    dp_13
        dp_5
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_457), .d2(_464), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_466[191:128]), .q2(_466[127:64]), .q1(_466[63:0]) );
    assign _469 = _466[63:0];
    assign data_19 = _469;
    assign address_22 = PHASE_4 ? _164 : _68;
    assign _533 = ~ PHASE_4;
    assign _532 = _70[6:6];
    assign read_enable_18 = _532 & _533;
    always @(posedge _84) begin
        if (_82)
            _503 <= _502;
        else
            _503 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _506 <= _505;
        else
            _506 <= _503;
    end
    always @(posedge _84) begin
        if (_82)
            _509 <= _508;
        else
            _509 <= _506;
    end
    always @(posedge _84) begin
        if (_82)
            _512 <= _511;
        else
            _512 <= _509;
    end
    always @(posedge _84) begin
        if (_82)
            _515 <= _514;
        else
            _515 <= _512;
    end
    always @(posedge _84) begin
        if (_82)
            _518 <= _517;
        else
            _518 <= _515;
    end
    always @(posedge _84) begin
        if (_82)
            _521 <= _520;
        else
            _521 <= _518;
    end
    always @(posedge _84) begin
        if (_82)
            _524 <= _523;
        else
            _524 <= _521;
    end
    always @(posedge _84) begin
        if (_82)
            _527 <= _526;
        else
            _527 <= _524;
    end
    assign _528 = ~ _527;
    always @(posedge _84) begin
        if (_82)
            _476 <= _475;
        else
            _476 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _479 <= _478;
        else
            _479 <= _476;
    end
    always @(posedge _84) begin
        if (_82)
            _482 <= _481;
        else
            _482 <= _479;
    end
    always @(posedge _84) begin
        if (_82)
            _485 <= _484;
        else
            _485 <= _482;
    end
    always @(posedge _84) begin
        if (_82)
            _488 <= _487;
        else
            _488 <= _485;
    end
    always @(posedge _84) begin
        if (_82)
            _491 <= _490;
        else
            _491 <= _488;
    end
    always @(posedge _84) begin
        if (_82)
            _494 <= _493;
        else
            _494 <= _491;
    end
    always @(posedge _84) begin
        if (_82)
            _497 <= _496;
        else
            _497 <= _494;
    end
    always @(posedge _84) begin
        if (_82)
            _500 <= _499;
        else
            _500 <= _497;
    end
    assign _529 = _500 & _528;
    assign _530 = _129 & _529;
    assign write_enable_22 = _530 & PHASE_4;
    assign _535 = write_enable_22 | read_enable_18;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_10
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_535), .regcea(vdd), .wea(write_enable_22), .addra(address_22), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_13), .regceb(vdd), .web(write_enable_13), .addrb(address_13), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_542[131:131]), .sbiterrb(_542[130:130]), .doutb(_542[129:66]), .dbiterra(_542[65:65]), .sbiterra(_542[64:64]), .douta(_542[63:0]) );
    assign _543 = _542[63:0];
    assign _473 = ~ PHASE_4;
    assign _15 = _473;
    always @(posedge _84) begin
        if (_82)
            PHASE_4 <= _471;
        else
            if (_72)
                PHASE_4 <= _15;
    end
    assign _555 = PHASE_4 ? _554 : _543;
    assign address_23 = _728 ? _199 : _723;
    assign write_enable_23 = _721 & _728;
    assign address_24 = _728 ? _164 : _68;
    assign _730 = ~ _728;
    assign read_enable_19 = _716 & _730;
    assign _728 = ~ PHASE_7;
    assign write_enable_24 = _714 & _728;
    assign _732 = write_enable_24 | read_enable_19;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_11
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_732), .regcea(vdd), .wea(write_enable_24), .addra(address_24), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_23), .regceb(vdd), .web(write_enable_23), .addrb(address_23), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_737[131:131]), .sbiterrb(_737[130:130]), .doutb(_737[129:66]), .dbiterra(_737[65:65]), .sbiterra(_737[64:64]), .douta(_737[63:0]) );
    assign _738 = _737[63:0];
    assign address_25 = PHASE_7 ? _199 : _723;
    assign _721 = _129 & _684;
    assign write_enable_25 = _721 & PHASE_7;
    assign _646 = _638[129:66];
    assign _645 = _625[129:66];
    assign _647 = PHASE_5 ? _646 : _645;
    assign _643 = _595[129:66];
    assign _642 = _581[129:66];
    assign q1_1 = PHASE_6 ? _643 : _642;
    assign _648 = _562 ? _647 : q1_1;
    assign address_26 = _627 ? _621 : _620;
    assign _633 = ~ _627;
    assign read_enable_20 = _102 & _633;
    assign address_27 = _627 ? _60 : _609;
    assign _629 = ~ _627;
    assign read_enable_21 = _102 & _629;
    assign _627 = ~ PHASE_5;
    assign write_enable_27 = _598 & _627;
    assign _631 = write_enable_27 | read_enable_21;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_12
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_631), .regcea(vdd), .wea(write_enable_27), .addra(address_27), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_20), .regceb(vdd), .web(write_enable_26), .addrb(address_26), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_638[131:131]), .sbiterrb(_638[130:130]), .doutb(_638[129:66]), .dbiterra(_638[65:65]), .sbiterra(_638[64:64]), .douta(_638[63:0]) );
    assign _639 = _638[63:0];
    assign _619 = _172[5:5];
    assign _618 = _172[4:4];
    assign _617 = _172[3:3];
    assign _616 = _172[2:2];
    assign _615 = _172[1:1];
    assign _614 = _172[0:0];
    assign _620 = { _614, _615, _616, _617, _618, _619 };
    assign address_28 = PHASE_5 ? _621 : _620;
    assign _611 = ~ PHASE_5;
    assign read_enable_22 = _102 & _611;
    assign data_25 = wr_d5;
    assign _608 = _137[5:5];
    assign _607 = _137[4:4];
    assign _606 = _137[3:3];
    assign _605 = _137[2:2];
    assign _604 = _137[1:1];
    assign _603 = _137[0:0];
    assign _609 = { _603, _604, _605, _606, _607, _608 };
    assign address_29 = PHASE_5 ? _60 : _609;
    assign _600 = ~ PHASE_5;
    assign read_enable_23 = _102 & _600;
    assign _598 = _62[5:5];
    assign write_enable_29 = _598 & PHASE_5;
    assign _602 = write_enable_29 | read_enable_23;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_13
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_602), .regcea(vdd), .wea(write_enable_29), .addra(address_29), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_22), .regceb(vdd), .web(write_enable_28), .addrb(address_28), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_625[131:131]), .sbiterrb(_625[130:130]), .doutb(_625[129:66]), .dbiterra(_625[65:65]), .sbiterra(_625[64:64]), .douta(_625[63:0]) );
    assign _626 = _625[63:0];
    assign _559 = ~ PHASE_5;
    assign _19 = _559;
    always @(posedge _84) begin
        if (_82)
            PHASE_5 <= _557;
        else
            if (_72)
                PHASE_5 <= _19;
    end
    assign _640 = PHASE_5 ? _639 : _626;
    assign address_30 = _583 ? _199 : _172;
    assign _590 = ~ _583;
    assign read_enable_24 = _102 & _590;
    assign write_enable_30 = _574 & _583;
    assign _592 = write_enable_30 | read_enable_24;
    assign address_31 = _583 ? _164 : _137;
    assign _585 = ~ _583;
    assign read_enable_25 = _102 & _585;
    assign _583 = ~ PHASE_6;
    assign write_enable_31 = _567 & _583;
    assign _587 = write_enable_31 | read_enable_25;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_14
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_587), .regcea(vdd), .wea(write_enable_31), .addra(address_31), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_592), .regceb(vdd), .web(write_enable_30), .addrb(address_30), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_595[131:131]), .sbiterrb(_595[130:130]), .doutb(_595[129:66]), .dbiterra(_595[65:65]), .sbiterra(_595[64:64]), .douta(_595[63:0]) );
    assign _596 = _595[63:0];
    assign _651 = _650[127:64];
    assign data_27 = _651;
    assign address_32 = PHASE_6 ? _199 : _172;
    assign _576 = ~ PHASE_6;
    assign read_enable_26 = _102 & _576;
    assign _573 = ~ _130;
    assign _574 = _129 & _573;
    assign write_enable_32 = _574 & PHASE_6;
    assign _578 = write_enable_32 | read_enable_26;
    assign address_33 = PHASE_6 ? _164 : _137;
    assign _569 = ~ PHASE_6;
    assign read_enable_27 = _102 & _569;
    assign _566 = ~ _130;
    assign _567 = _129 & _566;
    assign write_enable_33 = _567 & PHASE_6;
    assign _571 = write_enable_33 | read_enable_27;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_15
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_571), .regcea(vdd), .wea(write_enable_33), .addra(address_33), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_578), .regceb(vdd), .web(write_enable_32), .addrb(address_32), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_581[131:131]), .sbiterrb(_581[130:130]), .doutb(_581[129:66]), .dbiterra(_581[65:65]), .sbiterra(_581[64:64]), .douta(_581[63:0]) );
    assign _582 = _581[63:0];
    assign _652 = ~ PHASE_6;
    assign _21 = _652;
    always @(posedge _84) begin
        if (_82)
            PHASE_6 <= _564;
        else
            if (_99)
                PHASE_6 <= _21;
    end
    assign q0_1 = PHASE_6 ? _596 : _582;
    always @(posedge _84) begin
        if (_82)
            _562 <= _561;
        else
            _562 <= _92;
    end
    assign _641 = _562 ? _640 : q0_1;
    dp_12
        dp_4
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_641), .d2(_648), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_650[191:128]), .q2(_650[127:64]), .q1(_650[63:0]) );
    assign _653 = _650[63:0];
    assign data_31 = _653;
    assign address_34 = PHASE_7 ? _164 : _68;
    assign _717 = ~ PHASE_7;
    assign _716 = _70[5:5];
    assign read_enable_28 = _716 & _717;
    always @(posedge _84) begin
        if (_82)
            _687 <= _686;
        else
            _687 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _690 <= _689;
        else
            _690 <= _687;
    end
    always @(posedge _84) begin
        if (_82)
            _693 <= _692;
        else
            _693 <= _690;
    end
    always @(posedge _84) begin
        if (_82)
            _696 <= _695;
        else
            _696 <= _693;
    end
    always @(posedge _84) begin
        if (_82)
            _699 <= _698;
        else
            _699 <= _696;
    end
    always @(posedge _84) begin
        if (_82)
            _702 <= _701;
        else
            _702 <= _699;
    end
    always @(posedge _84) begin
        if (_82)
            _705 <= _704;
        else
            _705 <= _702;
    end
    always @(posedge _84) begin
        if (_82)
            _708 <= _707;
        else
            _708 <= _705;
    end
    always @(posedge _84) begin
        if (_82)
            _711 <= _710;
        else
            _711 <= _708;
    end
    assign _712 = ~ _711;
    always @(posedge _84) begin
        if (_82)
            _660 <= _659;
        else
            _660 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _663 <= _662;
        else
            _663 <= _660;
    end
    always @(posedge _84) begin
        if (_82)
            _666 <= _665;
        else
            _666 <= _663;
    end
    always @(posedge _84) begin
        if (_82)
            _669 <= _668;
        else
            _669 <= _666;
    end
    always @(posedge _84) begin
        if (_82)
            _672 <= _671;
        else
            _672 <= _669;
    end
    always @(posedge _84) begin
        if (_82)
            _675 <= _674;
        else
            _675 <= _672;
    end
    always @(posedge _84) begin
        if (_82)
            _678 <= _677;
        else
            _678 <= _675;
    end
    always @(posedge _84) begin
        if (_82)
            _681 <= _680;
        else
            _681 <= _678;
    end
    always @(posedge _84) begin
        if (_82)
            _684 <= _683;
        else
            _684 <= _681;
    end
    assign _713 = _684 & _712;
    assign _714 = _129 & _713;
    assign write_enable_34 = _714 & PHASE_7;
    assign _719 = write_enable_34 | read_enable_28;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_16
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_719), .regcea(vdd), .wea(write_enable_34), .addra(address_34), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_25), .regceb(vdd), .web(write_enable_25), .addrb(address_25), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_726[131:131]), .sbiterrb(_726[130:130]), .doutb(_726[129:66]), .dbiterra(_726[65:65]), .sbiterra(_726[64:64]), .douta(_726[63:0]) );
    assign _727 = _726[63:0];
    assign _657 = ~ PHASE_7;
    assign _23 = _657;
    always @(posedge _84) begin
        if (_82)
            PHASE_7 <= _655;
        else
            if (_72)
                PHASE_7 <= _23;
    end
    assign _739 = PHASE_7 ? _738 : _727;
    assign address_35 = _912 ? _199 : _907;
    assign write_enable_35 = _905 & _912;
    assign address_36 = _912 ? _164 : _68;
    assign _914 = ~ _912;
    assign read_enable_29 = _900 & _914;
    assign _912 = ~ PHASE_10;
    assign write_enable_36 = _898 & _912;
    assign _916 = write_enable_36 | read_enable_29;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_17
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_916), .regcea(vdd), .wea(write_enable_36), .addra(address_36), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_35), .regceb(vdd), .web(write_enable_35), .addrb(address_35), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_921[131:131]), .sbiterrb(_921[130:130]), .doutb(_921[129:66]), .dbiterra(_921[65:65]), .sbiterra(_921[64:64]), .douta(_921[63:0]) );
    assign _922 = _921[63:0];
    assign address_37 = PHASE_10 ? _199 : _907;
    assign _905 = _129 & _868;
    assign write_enable_37 = _905 & PHASE_10;
    assign _830 = _822[129:66];
    assign _829 = _809[129:66];
    assign _831 = PHASE_8 ? _830 : _829;
    assign _827 = _779[129:66];
    assign _826 = _765[129:66];
    assign q1_2 = PHASE_9 ? _827 : _826;
    assign _832 = _746 ? _831 : q1_2;
    assign address_38 = _811 ? _805 : _804;
    assign _817 = ~ _811;
    assign read_enable_30 = _102 & _817;
    assign address_39 = _811 ? _60 : _793;
    assign _813 = ~ _811;
    assign read_enable_31 = _102 & _813;
    assign _811 = ~ PHASE_8;
    assign write_enable_39 = _782 & _811;
    assign _815 = write_enable_39 | read_enable_31;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_18
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_815), .regcea(vdd), .wea(write_enable_39), .addra(address_39), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_30), .regceb(vdd), .web(write_enable_38), .addrb(address_38), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_822[131:131]), .sbiterrb(_822[130:130]), .doutb(_822[129:66]), .dbiterra(_822[65:65]), .sbiterra(_822[64:64]), .douta(_822[63:0]) );
    assign _823 = _822[63:0];
    assign _803 = _172[5:5];
    assign _802 = _172[4:4];
    assign _801 = _172[3:3];
    assign _800 = _172[2:2];
    assign _799 = _172[1:1];
    assign _798 = _172[0:0];
    assign _804 = { _798, _799, _800, _801, _802, _803 };
    assign address_40 = PHASE_8 ? _805 : _804;
    assign _795 = ~ PHASE_8;
    assign read_enable_32 = _102 & _795;
    assign data_37 = wr_d4;
    assign _792 = _137[5:5];
    assign _791 = _137[4:4];
    assign _790 = _137[3:3];
    assign _789 = _137[2:2];
    assign _788 = _137[1:1];
    assign _787 = _137[0:0];
    assign _793 = { _787, _788, _789, _790, _791, _792 };
    assign address_41 = PHASE_8 ? _60 : _793;
    assign _784 = ~ PHASE_8;
    assign read_enable_33 = _102 & _784;
    assign _782 = _62[4:4];
    assign write_enable_41 = _782 & PHASE_8;
    assign _786 = write_enable_41 | read_enable_33;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_19
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_786), .regcea(vdd), .wea(write_enable_41), .addra(address_41), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_32), .regceb(vdd), .web(write_enable_40), .addrb(address_40), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_809[131:131]), .sbiterrb(_809[130:130]), .doutb(_809[129:66]), .dbiterra(_809[65:65]), .sbiterra(_809[64:64]), .douta(_809[63:0]) );
    assign _810 = _809[63:0];
    assign _743 = ~ PHASE_8;
    assign _27 = _743;
    always @(posedge _84) begin
        if (_82)
            PHASE_8 <= _741;
        else
            if (_72)
                PHASE_8 <= _27;
    end
    assign _824 = PHASE_8 ? _823 : _810;
    assign address_42 = _767 ? _199 : _172;
    assign _774 = ~ _767;
    assign read_enable_34 = _102 & _774;
    assign write_enable_42 = _758 & _767;
    assign _776 = write_enable_42 | read_enable_34;
    assign address_43 = _767 ? _164 : _137;
    assign _769 = ~ _767;
    assign read_enable_35 = _102 & _769;
    assign _767 = ~ PHASE_9;
    assign write_enable_43 = _751 & _767;
    assign _771 = write_enable_43 | read_enable_35;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_20
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_771), .regcea(vdd), .wea(write_enable_43), .addra(address_43), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_776), .regceb(vdd), .web(write_enable_42), .addrb(address_42), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_779[131:131]), .sbiterrb(_779[130:130]), .doutb(_779[129:66]), .dbiterra(_779[65:65]), .sbiterra(_779[64:64]), .douta(_779[63:0]) );
    assign _780 = _779[63:0];
    assign _835 = _834[127:64];
    assign data_39 = _835;
    assign address_44 = PHASE_9 ? _199 : _172;
    assign _760 = ~ PHASE_9;
    assign read_enable_36 = _102 & _760;
    assign _757 = ~ _130;
    assign _758 = _129 & _757;
    assign write_enable_44 = _758 & PHASE_9;
    assign _762 = write_enable_44 | read_enable_36;
    assign address_45 = PHASE_9 ? _164 : _137;
    assign _753 = ~ PHASE_9;
    assign read_enable_37 = _102 & _753;
    assign _750 = ~ _130;
    assign _751 = _129 & _750;
    assign write_enable_45 = _751 & PHASE_9;
    assign _755 = write_enable_45 | read_enable_37;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_21
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_755), .regcea(vdd), .wea(write_enable_45), .addra(address_45), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_762), .regceb(vdd), .web(write_enable_44), .addrb(address_44), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_765[131:131]), .sbiterrb(_765[130:130]), .doutb(_765[129:66]), .dbiterra(_765[65:65]), .sbiterra(_765[64:64]), .douta(_765[63:0]) );
    assign _766 = _765[63:0];
    assign _836 = ~ PHASE_9;
    assign _29 = _836;
    always @(posedge _84) begin
        if (_82)
            PHASE_9 <= _748;
        else
            if (_99)
                PHASE_9 <= _29;
    end
    assign q0_2 = PHASE_9 ? _780 : _766;
    always @(posedge _84) begin
        if (_82)
            _746 <= _745;
        else
            _746 <= _92;
    end
    assign _825 = _746 ? _824 : q0_2;
    dp_11
        dp_3
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_825), .d2(_832), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_834[191:128]), .q2(_834[127:64]), .q1(_834[63:0]) );
    assign _837 = _834[63:0];
    assign data_43 = _837;
    assign address_46 = PHASE_10 ? _164 : _68;
    assign _901 = ~ PHASE_10;
    assign _900 = _70[4:4];
    assign read_enable_38 = _900 & _901;
    always @(posedge _84) begin
        if (_82)
            _871 <= _870;
        else
            _871 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _874 <= _873;
        else
            _874 <= _871;
    end
    always @(posedge _84) begin
        if (_82)
            _877 <= _876;
        else
            _877 <= _874;
    end
    always @(posedge _84) begin
        if (_82)
            _880 <= _879;
        else
            _880 <= _877;
    end
    always @(posedge _84) begin
        if (_82)
            _883 <= _882;
        else
            _883 <= _880;
    end
    always @(posedge _84) begin
        if (_82)
            _886 <= _885;
        else
            _886 <= _883;
    end
    always @(posedge _84) begin
        if (_82)
            _889 <= _888;
        else
            _889 <= _886;
    end
    always @(posedge _84) begin
        if (_82)
            _892 <= _891;
        else
            _892 <= _889;
    end
    always @(posedge _84) begin
        if (_82)
            _895 <= _894;
        else
            _895 <= _892;
    end
    assign _896 = ~ _895;
    always @(posedge _84) begin
        if (_82)
            _844 <= _843;
        else
            _844 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _847 <= _846;
        else
            _847 <= _844;
    end
    always @(posedge _84) begin
        if (_82)
            _850 <= _849;
        else
            _850 <= _847;
    end
    always @(posedge _84) begin
        if (_82)
            _853 <= _852;
        else
            _853 <= _850;
    end
    always @(posedge _84) begin
        if (_82)
            _856 <= _855;
        else
            _856 <= _853;
    end
    always @(posedge _84) begin
        if (_82)
            _859 <= _858;
        else
            _859 <= _856;
    end
    always @(posedge _84) begin
        if (_82)
            _862 <= _861;
        else
            _862 <= _859;
    end
    always @(posedge _84) begin
        if (_82)
            _865 <= _864;
        else
            _865 <= _862;
    end
    always @(posedge _84) begin
        if (_82)
            _868 <= _867;
        else
            _868 <= _865;
    end
    assign _897 = _868 & _896;
    assign _898 = _129 & _897;
    assign write_enable_46 = _898 & PHASE_10;
    assign _903 = write_enable_46 | read_enable_38;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_22
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_903), .regcea(vdd), .wea(write_enable_46), .addra(address_46), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_37), .regceb(vdd), .web(write_enable_37), .addrb(address_37), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_910[131:131]), .sbiterrb(_910[130:130]), .doutb(_910[129:66]), .dbiterra(_910[65:65]), .sbiterra(_910[64:64]), .douta(_910[63:0]) );
    assign _911 = _910[63:0];
    assign _841 = ~ PHASE_10;
    assign _31 = _841;
    always @(posedge _84) begin
        if (_82)
            PHASE_10 <= _839;
        else
            if (_72)
                PHASE_10 <= _31;
    end
    assign _923 = PHASE_10 ? _922 : _911;
    assign address_47 = _1096 ? _199 : _1091;
    assign write_enable_47 = _1089 & _1096;
    assign address_48 = _1096 ? _164 : _68;
    assign _1098 = ~ _1096;
    assign read_enable_39 = _1084 & _1098;
    assign _1096 = ~ PHASE_13;
    assign write_enable_48 = _1082 & _1096;
    assign _1100 = write_enable_48 | read_enable_39;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_23
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1100), .regcea(vdd), .wea(write_enable_48), .addra(address_48), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_47), .regceb(vdd), .web(write_enable_47), .addrb(address_47), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1105[131:131]), .sbiterrb(_1105[130:130]), .doutb(_1105[129:66]), .dbiterra(_1105[65:65]), .sbiterra(_1105[64:64]), .douta(_1105[63:0]) );
    assign _1106 = _1105[63:0];
    assign address_49 = PHASE_13 ? _199 : _1091;
    assign _1089 = _129 & _1052;
    assign write_enable_49 = _1089 & PHASE_13;
    assign _1014 = _1006[129:66];
    assign _1013 = _993[129:66];
    assign _1015 = PHASE_11 ? _1014 : _1013;
    assign _1011 = _963[129:66];
    assign _1010 = _949[129:66];
    assign q1_3 = PHASE_12 ? _1011 : _1010;
    assign _1016 = _930 ? _1015 : q1_3;
    assign address_50 = _995 ? _989 : _988;
    assign _1001 = ~ _995;
    assign read_enable_40 = _102 & _1001;
    assign address_51 = _995 ? _60 : _977;
    assign _997 = ~ _995;
    assign read_enable_41 = _102 & _997;
    assign _995 = ~ PHASE_11;
    assign write_enable_51 = _966 & _995;
    assign _999 = write_enable_51 | read_enable_41;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_24
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_999), .regcea(vdd), .wea(write_enable_51), .addra(address_51), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_40), .regceb(vdd), .web(write_enable_50), .addrb(address_50), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1006[131:131]), .sbiterrb(_1006[130:130]), .doutb(_1006[129:66]), .dbiterra(_1006[65:65]), .sbiterra(_1006[64:64]), .douta(_1006[63:0]) );
    assign _1007 = _1006[63:0];
    assign _987 = _172[5:5];
    assign _986 = _172[4:4];
    assign _985 = _172[3:3];
    assign _984 = _172[2:2];
    assign _983 = _172[1:1];
    assign _982 = _172[0:0];
    assign _988 = { _982, _983, _984, _985, _986, _987 };
    assign address_52 = PHASE_11 ? _989 : _988;
    assign _979 = ~ PHASE_11;
    assign read_enable_42 = _102 & _979;
    assign data_49 = wr_d3;
    assign _976 = _137[5:5];
    assign _975 = _137[4:4];
    assign _974 = _137[3:3];
    assign _973 = _137[2:2];
    assign _972 = _137[1:1];
    assign _971 = _137[0:0];
    assign _977 = { _971, _972, _973, _974, _975, _976 };
    assign address_53 = PHASE_11 ? _60 : _977;
    assign _968 = ~ PHASE_11;
    assign read_enable_43 = _102 & _968;
    assign _966 = _62[3:3];
    assign write_enable_53 = _966 & PHASE_11;
    assign _970 = write_enable_53 | read_enable_43;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_25
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_970), .regcea(vdd), .wea(write_enable_53), .addra(address_53), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_42), .regceb(vdd), .web(write_enable_52), .addrb(address_52), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_993[131:131]), .sbiterrb(_993[130:130]), .doutb(_993[129:66]), .dbiterra(_993[65:65]), .sbiterra(_993[64:64]), .douta(_993[63:0]) );
    assign _994 = _993[63:0];
    assign _927 = ~ PHASE_11;
    assign _35 = _927;
    always @(posedge _84) begin
        if (_82)
            PHASE_11 <= _925;
        else
            if (_72)
                PHASE_11 <= _35;
    end
    assign _1008 = PHASE_11 ? _1007 : _994;
    assign address_54 = _951 ? _199 : _172;
    assign _958 = ~ _951;
    assign read_enable_44 = _102 & _958;
    assign write_enable_54 = _942 & _951;
    assign _960 = write_enable_54 | read_enable_44;
    assign address_55 = _951 ? _164 : _137;
    assign _953 = ~ _951;
    assign read_enable_45 = _102 & _953;
    assign _951 = ~ PHASE_12;
    assign write_enable_55 = _935 & _951;
    assign _955 = write_enable_55 | read_enable_45;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_26
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_955), .regcea(vdd), .wea(write_enable_55), .addra(address_55), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_960), .regceb(vdd), .web(write_enable_54), .addrb(address_54), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_963[131:131]), .sbiterrb(_963[130:130]), .doutb(_963[129:66]), .dbiterra(_963[65:65]), .sbiterra(_963[64:64]), .douta(_963[63:0]) );
    assign _964 = _963[63:0];
    assign _1019 = _1018[127:64];
    assign data_51 = _1019;
    assign address_56 = PHASE_12 ? _199 : _172;
    assign _944 = ~ PHASE_12;
    assign read_enable_46 = _102 & _944;
    assign _941 = ~ _130;
    assign _942 = _129 & _941;
    assign write_enable_56 = _942 & PHASE_12;
    assign _946 = write_enable_56 | read_enable_46;
    assign address_57 = PHASE_12 ? _164 : _137;
    assign _937 = ~ PHASE_12;
    assign read_enable_47 = _102 & _937;
    assign _934 = ~ _130;
    assign _935 = _129 & _934;
    assign write_enable_57 = _935 & PHASE_12;
    assign _939 = write_enable_57 | read_enable_47;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_27
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_939), .regcea(vdd), .wea(write_enable_57), .addra(address_57), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_946), .regceb(vdd), .web(write_enable_56), .addrb(address_56), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_949[131:131]), .sbiterrb(_949[130:130]), .doutb(_949[129:66]), .dbiterra(_949[65:65]), .sbiterra(_949[64:64]), .douta(_949[63:0]) );
    assign _950 = _949[63:0];
    assign _1020 = ~ PHASE_12;
    assign _37 = _1020;
    always @(posedge _84) begin
        if (_82)
            PHASE_12 <= _932;
        else
            if (_99)
                PHASE_12 <= _37;
    end
    assign q0_3 = PHASE_12 ? _964 : _950;
    always @(posedge _84) begin
        if (_82)
            _930 <= _929;
        else
            _930 <= _92;
    end
    assign _1009 = _930 ? _1008 : q0_3;
    dp_10
        dp_2
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1009), .d2(_1016), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_1018[191:128]), .q2(_1018[127:64]), .q1(_1018[63:0]) );
    assign _1021 = _1018[63:0];
    assign data_55 = _1021;
    assign address_58 = PHASE_13 ? _164 : _68;
    assign _1085 = ~ PHASE_13;
    assign _1084 = _70[3:3];
    assign read_enable_48 = _1084 & _1085;
    always @(posedge _84) begin
        if (_82)
            _1055 <= _1054;
        else
            _1055 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _1058 <= _1057;
        else
            _1058 <= _1055;
    end
    always @(posedge _84) begin
        if (_82)
            _1061 <= _1060;
        else
            _1061 <= _1058;
    end
    always @(posedge _84) begin
        if (_82)
            _1064 <= _1063;
        else
            _1064 <= _1061;
    end
    always @(posedge _84) begin
        if (_82)
            _1067 <= _1066;
        else
            _1067 <= _1064;
    end
    always @(posedge _84) begin
        if (_82)
            _1070 <= _1069;
        else
            _1070 <= _1067;
    end
    always @(posedge _84) begin
        if (_82)
            _1073 <= _1072;
        else
            _1073 <= _1070;
    end
    always @(posedge _84) begin
        if (_82)
            _1076 <= _1075;
        else
            _1076 <= _1073;
    end
    always @(posedge _84) begin
        if (_82)
            _1079 <= _1078;
        else
            _1079 <= _1076;
    end
    assign _1080 = ~ _1079;
    always @(posedge _84) begin
        if (_82)
            _1028 <= _1027;
        else
            _1028 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1031 <= _1030;
        else
            _1031 <= _1028;
    end
    always @(posedge _84) begin
        if (_82)
            _1034 <= _1033;
        else
            _1034 <= _1031;
    end
    always @(posedge _84) begin
        if (_82)
            _1037 <= _1036;
        else
            _1037 <= _1034;
    end
    always @(posedge _84) begin
        if (_82)
            _1040 <= _1039;
        else
            _1040 <= _1037;
    end
    always @(posedge _84) begin
        if (_82)
            _1043 <= _1042;
        else
            _1043 <= _1040;
    end
    always @(posedge _84) begin
        if (_82)
            _1046 <= _1045;
        else
            _1046 <= _1043;
    end
    always @(posedge _84) begin
        if (_82)
            _1049 <= _1048;
        else
            _1049 <= _1046;
    end
    always @(posedge _84) begin
        if (_82)
            _1052 <= _1051;
        else
            _1052 <= _1049;
    end
    assign _1081 = _1052 & _1080;
    assign _1082 = _129 & _1081;
    assign write_enable_58 = _1082 & PHASE_13;
    assign _1087 = write_enable_58 | read_enable_48;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_28
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1087), .regcea(vdd), .wea(write_enable_58), .addra(address_58), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_49), .regceb(vdd), .web(write_enable_49), .addrb(address_49), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1094[131:131]), .sbiterrb(_1094[130:130]), .doutb(_1094[129:66]), .dbiterra(_1094[65:65]), .sbiterra(_1094[64:64]), .douta(_1094[63:0]) );
    assign _1095 = _1094[63:0];
    assign _1025 = ~ PHASE_13;
    assign _39 = _1025;
    always @(posedge _84) begin
        if (_82)
            PHASE_13 <= _1023;
        else
            if (_72)
                PHASE_13 <= _39;
    end
    assign _1107 = PHASE_13 ? _1106 : _1095;
    assign address_59 = _1280 ? _199 : _1275;
    assign write_enable_59 = _1273 & _1280;
    assign address_60 = _1280 ? _164 : _68;
    assign _1282 = ~ _1280;
    assign read_enable_49 = _1268 & _1282;
    assign _1280 = ~ PHASE_16;
    assign write_enable_60 = _1266 & _1280;
    assign _1284 = write_enable_60 | read_enable_49;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_29
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1284), .regcea(vdd), .wea(write_enable_60), .addra(address_60), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_59), .regceb(vdd), .web(write_enable_59), .addrb(address_59), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1289[131:131]), .sbiterrb(_1289[130:130]), .doutb(_1289[129:66]), .dbiterra(_1289[65:65]), .sbiterra(_1289[64:64]), .douta(_1289[63:0]) );
    assign _1290 = _1289[63:0];
    assign address_61 = PHASE_16 ? _199 : _1275;
    assign _1273 = _129 & _1236;
    assign write_enable_61 = _1273 & PHASE_16;
    assign _1198 = _1190[129:66];
    assign _1197 = _1177[129:66];
    assign _1199 = PHASE_14 ? _1198 : _1197;
    assign _1195 = _1147[129:66];
    assign _1194 = _1133[129:66];
    assign q1_4 = PHASE_15 ? _1195 : _1194;
    assign _1200 = _1114 ? _1199 : q1_4;
    assign address_62 = _1179 ? _1173 : _1172;
    assign _1185 = ~ _1179;
    assign read_enable_50 = _102 & _1185;
    assign address_63 = _1179 ? _60 : _1161;
    assign _1181 = ~ _1179;
    assign read_enable_51 = _102 & _1181;
    assign _1179 = ~ PHASE_14;
    assign write_enable_63 = _1150 & _1179;
    assign _1183 = write_enable_63 | read_enable_51;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_30
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1183), .regcea(vdd), .wea(write_enable_63), .addra(address_63), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_50), .regceb(vdd), .web(write_enable_62), .addrb(address_62), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1190[131:131]), .sbiterrb(_1190[130:130]), .doutb(_1190[129:66]), .dbiterra(_1190[65:65]), .sbiterra(_1190[64:64]), .douta(_1190[63:0]) );
    assign _1191 = _1190[63:0];
    assign _1171 = _172[5:5];
    assign _1170 = _172[4:4];
    assign _1169 = _172[3:3];
    assign _1168 = _172[2:2];
    assign _1167 = _172[1:1];
    assign _1166 = _172[0:0];
    assign _1172 = { _1166, _1167, _1168, _1169, _1170, _1171 };
    assign address_64 = PHASE_14 ? _1173 : _1172;
    assign _1163 = ~ PHASE_14;
    assign read_enable_52 = _102 & _1163;
    assign data_61 = wr_d2;
    assign _1160 = _137[5:5];
    assign _1159 = _137[4:4];
    assign _1158 = _137[3:3];
    assign _1157 = _137[2:2];
    assign _1156 = _137[1:1];
    assign _1155 = _137[0:0];
    assign _1161 = { _1155, _1156, _1157, _1158, _1159, _1160 };
    assign address_65 = PHASE_14 ? _60 : _1161;
    assign _1152 = ~ PHASE_14;
    assign read_enable_53 = _102 & _1152;
    assign _1150 = _62[2:2];
    assign write_enable_65 = _1150 & PHASE_14;
    assign _1154 = write_enable_65 | read_enable_53;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_31
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1154), .regcea(vdd), .wea(write_enable_65), .addra(address_65), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_52), .regceb(vdd), .web(write_enable_64), .addrb(address_64), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1177[131:131]), .sbiterrb(_1177[130:130]), .doutb(_1177[129:66]), .dbiterra(_1177[65:65]), .sbiterra(_1177[64:64]), .douta(_1177[63:0]) );
    assign _1178 = _1177[63:0];
    assign _1111 = ~ PHASE_14;
    assign _43 = _1111;
    always @(posedge _84) begin
        if (_82)
            PHASE_14 <= _1109;
        else
            if (_72)
                PHASE_14 <= _43;
    end
    assign _1192 = PHASE_14 ? _1191 : _1178;
    assign address_66 = _1135 ? _199 : _172;
    assign _1142 = ~ _1135;
    assign read_enable_54 = _102 & _1142;
    assign write_enable_66 = _1126 & _1135;
    assign _1144 = write_enable_66 | read_enable_54;
    assign address_67 = _1135 ? _164 : _137;
    assign _1137 = ~ _1135;
    assign read_enable_55 = _102 & _1137;
    assign _1135 = ~ PHASE_15;
    assign write_enable_67 = _1119 & _1135;
    assign _1139 = write_enable_67 | read_enable_55;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_32
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1139), .regcea(vdd), .wea(write_enable_67), .addra(address_67), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1144), .regceb(vdd), .web(write_enable_66), .addrb(address_66), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1147[131:131]), .sbiterrb(_1147[130:130]), .doutb(_1147[129:66]), .dbiterra(_1147[65:65]), .sbiterra(_1147[64:64]), .douta(_1147[63:0]) );
    assign _1148 = _1147[63:0];
    assign _1203 = _1202[127:64];
    assign data_63 = _1203;
    assign address_68 = PHASE_15 ? _199 : _172;
    assign _1128 = ~ PHASE_15;
    assign read_enable_56 = _102 & _1128;
    assign _1125 = ~ _130;
    assign _1126 = _129 & _1125;
    assign write_enable_68 = _1126 & PHASE_15;
    assign _1130 = write_enable_68 | read_enable_56;
    assign address_69 = PHASE_15 ? _164 : _137;
    assign _1121 = ~ PHASE_15;
    assign read_enable_57 = _102 & _1121;
    assign _1118 = ~ _130;
    assign _1119 = _129 & _1118;
    assign write_enable_69 = _1119 & PHASE_15;
    assign _1123 = write_enable_69 | read_enable_57;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_33
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1123), .regcea(vdd), .wea(write_enable_69), .addra(address_69), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1130), .regceb(vdd), .web(write_enable_68), .addrb(address_68), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1133[131:131]), .sbiterrb(_1133[130:130]), .doutb(_1133[129:66]), .dbiterra(_1133[65:65]), .sbiterra(_1133[64:64]), .douta(_1133[63:0]) );
    assign _1134 = _1133[63:0];
    assign _1204 = ~ PHASE_15;
    assign _45 = _1204;
    always @(posedge _84) begin
        if (_82)
            PHASE_15 <= _1116;
        else
            if (_99)
                PHASE_15 <= _45;
    end
    assign q0_4 = PHASE_15 ? _1148 : _1134;
    always @(posedge _84) begin
        if (_82)
            _1114 <= _1113;
        else
            _1114 <= _92;
    end
    assign _1193 = _1114 ? _1192 : q0_4;
    dp_9
        dp_1
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1193), .d2(_1200), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_1202[191:128]), .q2(_1202[127:64]), .q1(_1202[63:0]) );
    assign _1205 = _1202[63:0];
    assign data_67 = _1205;
    assign address_70 = PHASE_16 ? _164 : _68;
    assign _1269 = ~ PHASE_16;
    assign _1268 = _70[2:2];
    assign read_enable_58 = _1268 & _1269;
    always @(posedge _84) begin
        if (_82)
            _1239 <= _1238;
        else
            _1239 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _1242 <= _1241;
        else
            _1242 <= _1239;
    end
    always @(posedge _84) begin
        if (_82)
            _1245 <= _1244;
        else
            _1245 <= _1242;
    end
    always @(posedge _84) begin
        if (_82)
            _1248 <= _1247;
        else
            _1248 <= _1245;
    end
    always @(posedge _84) begin
        if (_82)
            _1251 <= _1250;
        else
            _1251 <= _1248;
    end
    always @(posedge _84) begin
        if (_82)
            _1254 <= _1253;
        else
            _1254 <= _1251;
    end
    always @(posedge _84) begin
        if (_82)
            _1257 <= _1256;
        else
            _1257 <= _1254;
    end
    always @(posedge _84) begin
        if (_82)
            _1260 <= _1259;
        else
            _1260 <= _1257;
    end
    always @(posedge _84) begin
        if (_82)
            _1263 <= _1262;
        else
            _1263 <= _1260;
    end
    assign _1264 = ~ _1263;
    always @(posedge _84) begin
        if (_82)
            _1212 <= _1211;
        else
            _1212 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1215 <= _1214;
        else
            _1215 <= _1212;
    end
    always @(posedge _84) begin
        if (_82)
            _1218 <= _1217;
        else
            _1218 <= _1215;
    end
    always @(posedge _84) begin
        if (_82)
            _1221 <= _1220;
        else
            _1221 <= _1218;
    end
    always @(posedge _84) begin
        if (_82)
            _1224 <= _1223;
        else
            _1224 <= _1221;
    end
    always @(posedge _84) begin
        if (_82)
            _1227 <= _1226;
        else
            _1227 <= _1224;
    end
    always @(posedge _84) begin
        if (_82)
            _1230 <= _1229;
        else
            _1230 <= _1227;
    end
    always @(posedge _84) begin
        if (_82)
            _1233 <= _1232;
        else
            _1233 <= _1230;
    end
    always @(posedge _84) begin
        if (_82)
            _1236 <= _1235;
        else
            _1236 <= _1233;
    end
    assign _1265 = _1236 & _1264;
    assign _1266 = _129 & _1265;
    assign write_enable_70 = _1266 & PHASE_16;
    assign _1271 = write_enable_70 | read_enable_58;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_34
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1271), .regcea(vdd), .wea(write_enable_70), .addra(address_70), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_61), .regceb(vdd), .web(write_enable_61), .addrb(address_61), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1278[131:131]), .sbiterrb(_1278[130:130]), .doutb(_1278[129:66]), .dbiterra(_1278[65:65]), .sbiterra(_1278[64:64]), .douta(_1278[63:0]) );
    assign _1279 = _1278[63:0];
    assign _1209 = ~ PHASE_16;
    assign _47 = _1209;
    always @(posedge _84) begin
        if (_82)
            PHASE_16 <= _1207;
        else
            if (_72)
                PHASE_16 <= _47;
    end
    assign _1291 = PHASE_16 ? _1290 : _1279;
    assign address_71 = _1464 ? _199 : _1459;
    assign write_enable_71 = _1457 & _1464;
    assign address_72 = _1464 ? _164 : _68;
    assign _1466 = ~ _1464;
    assign read_enable_59 = _1452 & _1466;
    assign _1464 = ~ PHASE_19;
    assign write_enable_72 = _1450 & _1464;
    assign _1468 = write_enable_72 | read_enable_59;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_35
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1468), .regcea(vdd), .wea(write_enable_72), .addra(address_72), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_71), .regceb(vdd), .web(write_enable_71), .addrb(address_71), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1473[131:131]), .sbiterrb(_1473[130:130]), .doutb(_1473[129:66]), .dbiterra(_1473[65:65]), .sbiterra(_1473[64:64]), .douta(_1473[63:0]) );
    assign _1474 = _1473[63:0];
    assign address_73 = PHASE_19 ? _199 : _1459;
    assign _1457 = _129 & _1420;
    assign write_enable_73 = _1457 & PHASE_19;
    assign _1382 = _1374[129:66];
    assign _1381 = _1361[129:66];
    assign _1383 = PHASE_17 ? _1382 : _1381;
    assign _1379 = _1331[129:66];
    assign _1378 = _1317[129:66];
    assign q1_5 = PHASE_18 ? _1379 : _1378;
    assign _1384 = _1298 ? _1383 : q1_5;
    assign address_74 = _1363 ? _1357 : _1356;
    assign _1369 = ~ _1363;
    assign read_enable_60 = _102 & _1369;
    assign address_75 = _1363 ? _60 : _1345;
    assign _1365 = ~ _1363;
    assign read_enable_61 = _102 & _1365;
    assign _1363 = ~ PHASE_17;
    assign write_enable_75 = _1334 & _1363;
    assign _1367 = write_enable_75 | read_enable_61;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_36
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1367), .regcea(vdd), .wea(write_enable_75), .addra(address_75), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_60), .regceb(vdd), .web(write_enable_74), .addrb(address_74), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1374[131:131]), .sbiterrb(_1374[130:130]), .doutb(_1374[129:66]), .dbiterra(_1374[65:65]), .sbiterra(_1374[64:64]), .douta(_1374[63:0]) );
    assign _1375 = _1374[63:0];
    assign _1355 = _172[5:5];
    assign _1354 = _172[4:4];
    assign _1353 = _172[3:3];
    assign _1352 = _172[2:2];
    assign _1351 = _172[1:1];
    assign _1350 = _172[0:0];
    assign _1356 = { _1350, _1351, _1352, _1353, _1354, _1355 };
    assign address_76 = PHASE_17 ? _1357 : _1356;
    assign _1347 = ~ PHASE_17;
    assign read_enable_62 = _102 & _1347;
    assign data_73 = wr_d1;
    assign _1344 = _137[5:5];
    assign _1343 = _137[4:4];
    assign _1342 = _137[3:3];
    assign _1341 = _137[2:2];
    assign _1340 = _137[1:1];
    assign _1339 = _137[0:0];
    assign _1345 = { _1339, _1340, _1341, _1342, _1343, _1344 };
    assign address_77 = PHASE_17 ? _60 : _1345;
    assign _1336 = ~ PHASE_17;
    assign read_enable_63 = _102 & _1336;
    assign _1334 = _62[1:1];
    assign write_enable_77 = _1334 & PHASE_17;
    assign _1338 = write_enable_77 | read_enable_63;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_37
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1338), .regcea(vdd), .wea(write_enable_77), .addra(address_77), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_62), .regceb(vdd), .web(write_enable_76), .addrb(address_76), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1361[131:131]), .sbiterrb(_1361[130:130]), .doutb(_1361[129:66]), .dbiterra(_1361[65:65]), .sbiterra(_1361[64:64]), .douta(_1361[63:0]) );
    assign _1362 = _1361[63:0];
    assign _1295 = ~ PHASE_17;
    assign _51 = _1295;
    always @(posedge _84) begin
        if (_82)
            PHASE_17 <= _1293;
        else
            if (_72)
                PHASE_17 <= _51;
    end
    assign _1376 = PHASE_17 ? _1375 : _1362;
    assign address_78 = _1319 ? _199 : _172;
    assign _1326 = ~ _1319;
    assign read_enable_64 = _102 & _1326;
    assign write_enable_78 = _1310 & _1319;
    assign _1328 = write_enable_78 | read_enable_64;
    assign address_79 = _1319 ? _164 : _137;
    assign _1321 = ~ _1319;
    assign read_enable_65 = _102 & _1321;
    assign _1319 = ~ PHASE_18;
    assign write_enable_79 = _1303 & _1319;
    assign _1323 = write_enable_79 | read_enable_65;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_38
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1323), .regcea(vdd), .wea(write_enable_79), .addra(address_79), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1328), .regceb(vdd), .web(write_enable_78), .addrb(address_78), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1331[131:131]), .sbiterrb(_1331[130:130]), .doutb(_1331[129:66]), .dbiterra(_1331[65:65]), .sbiterra(_1331[64:64]), .douta(_1331[63:0]) );
    assign _1332 = _1331[63:0];
    assign _1387 = _1386[127:64];
    assign data_75 = _1387;
    assign address_80 = PHASE_18 ? _199 : _172;
    assign _1312 = ~ PHASE_18;
    assign read_enable_66 = _102 & _1312;
    assign _1309 = ~ _130;
    assign _1310 = _129 & _1309;
    assign write_enable_80 = _1310 & PHASE_18;
    assign _1314 = write_enable_80 | read_enable_66;
    assign address_81 = PHASE_18 ? _164 : _137;
    assign _1305 = ~ PHASE_18;
    assign read_enable_67 = _102 & _1305;
    assign _1302 = ~ _130;
    assign _1303 = _129 & _1302;
    assign write_enable_81 = _1303 & PHASE_18;
    assign _1307 = write_enable_81 | read_enable_67;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_39
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1307), .regcea(vdd), .wea(write_enable_81), .addra(address_81), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1314), .regceb(vdd), .web(write_enable_80), .addrb(address_80), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1317[131:131]), .sbiterrb(_1317[130:130]), .doutb(_1317[129:66]), .dbiterra(_1317[65:65]), .sbiterra(_1317[64:64]), .douta(_1317[63:0]) );
    assign _1318 = _1317[63:0];
    assign _1388 = ~ PHASE_18;
    assign _53 = _1388;
    always @(posedge _84) begin
        if (_82)
            PHASE_18 <= _1300;
        else
            if (_99)
                PHASE_18 <= _53;
    end
    assign q0_5 = PHASE_18 ? _1332 : _1318;
    always @(posedge _84) begin
        if (_82)
            _1298 <= _1297;
        else
            _1298 <= _92;
    end
    assign _1377 = _1298 ? _1376 : q0_5;
    dp_8
        dp_0
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1377), .d2(_1384), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_1386[191:128]), .q2(_1386[127:64]), .q1(_1386[63:0]) );
    assign _1389 = _1386[63:0];
    assign data_79 = _1389;
    assign address_82 = PHASE_19 ? _164 : _68;
    assign _1453 = ~ PHASE_19;
    assign _1452 = _70[1:1];
    assign read_enable_68 = _1452 & _1453;
    always @(posedge _84) begin
        if (_82)
            _1423 <= _1422;
        else
            _1423 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _1426 <= _1425;
        else
            _1426 <= _1423;
    end
    always @(posedge _84) begin
        if (_82)
            _1429 <= _1428;
        else
            _1429 <= _1426;
    end
    always @(posedge _84) begin
        if (_82)
            _1432 <= _1431;
        else
            _1432 <= _1429;
    end
    always @(posedge _84) begin
        if (_82)
            _1435 <= _1434;
        else
            _1435 <= _1432;
    end
    always @(posedge _84) begin
        if (_82)
            _1438 <= _1437;
        else
            _1438 <= _1435;
    end
    always @(posedge _84) begin
        if (_82)
            _1441 <= _1440;
        else
            _1441 <= _1438;
    end
    always @(posedge _84) begin
        if (_82)
            _1444 <= _1443;
        else
            _1444 <= _1441;
    end
    always @(posedge _84) begin
        if (_82)
            _1447 <= _1446;
        else
            _1447 <= _1444;
    end
    assign _1448 = ~ _1447;
    always @(posedge _84) begin
        if (_82)
            _1396 <= _1395;
        else
            _1396 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1399 <= _1398;
        else
            _1399 <= _1396;
    end
    always @(posedge _84) begin
        if (_82)
            _1402 <= _1401;
        else
            _1402 <= _1399;
    end
    always @(posedge _84) begin
        if (_82)
            _1405 <= _1404;
        else
            _1405 <= _1402;
    end
    always @(posedge _84) begin
        if (_82)
            _1408 <= _1407;
        else
            _1408 <= _1405;
    end
    always @(posedge _84) begin
        if (_82)
            _1411 <= _1410;
        else
            _1411 <= _1408;
    end
    always @(posedge _84) begin
        if (_82)
            _1414 <= _1413;
        else
            _1414 <= _1411;
    end
    always @(posedge _84) begin
        if (_82)
            _1417 <= _1416;
        else
            _1417 <= _1414;
    end
    always @(posedge _84) begin
        if (_82)
            _1420 <= _1419;
        else
            _1420 <= _1417;
    end
    assign _1449 = _1420 & _1448;
    assign _1450 = _129 & _1449;
    assign write_enable_82 = _1450 & PHASE_19;
    assign _1455 = write_enable_82 | read_enable_68;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_40
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1455), .regcea(vdd), .wea(write_enable_82), .addra(address_82), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_73), .regceb(vdd), .web(write_enable_73), .addrb(address_73), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1462[131:131]), .sbiterrb(_1462[130:130]), .doutb(_1462[129:66]), .dbiterra(_1462[65:65]), .sbiterra(_1462[64:64]), .douta(_1462[63:0]) );
    assign _1463 = _1462[63:0];
    assign _1393 = ~ PHASE_19;
    assign _55 = _1393;
    always @(posedge _84) begin
        if (_82)
            PHASE_19 <= _1391;
        else
            if (_72)
                PHASE_19 <= _55;
    end
    assign _1475 = PHASE_19 ? _1474 : _1463;
    assign address_83 = _1648 ? _199 : _1643;
    assign write_enable_83 = _1641 & _1648;
    assign address_84 = _1648 ? _164 : _68;
    assign _1650 = ~ _1648;
    assign read_enable_69 = _1636 & _1650;
    assign _1648 = ~ PHASE_22;
    assign write_enable_84 = _1634 & _1648;
    assign _1652 = write_enable_84 | read_enable_69;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_41
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1652), .regcea(vdd), .wea(write_enable_84), .addra(address_84), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_83), .regceb(vdd), .web(write_enable_83), .addrb(address_83), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1657[131:131]), .sbiterrb(_1657[130:130]), .doutb(_1657[129:66]), .dbiterra(_1657[65:65]), .sbiterra(_1657[64:64]), .douta(_1657[63:0]) );
    assign _1658 = _1657[63:0];
    assign address_85 = PHASE_22 ? _199 : _1643;
    assign _1641 = _129 & _1604;
    assign write_enable_85 = _1641 & PHASE_22;
    assign _280 = _91[490:487];
    assign _279 = _91[486:486];
    assign _277 = _91[482:482];
    assign _276 = _91[481:418];
    assign _275 = _91[417:354];
    assign _274 = _91[353:290];
    assign _273 = _91[289:226];
    assign _272 = _91[225:162];
    assign _271 = _91[161:98];
    assign _270 = _91[97:34];
    assign _1566 = _1558[129:66];
    assign _1565 = _1545[129:66];
    assign _1567 = PHASE_20 ? _1566 : _1565;
    assign _1563 = _1515[129:66];
    assign _1562 = _1501[129:66];
    assign q1_6 = PHASE_21 ? _1563 : _1562;
    assign _1568 = _1482 ? _1567 : q1_6;
    assign address_86 = _1547 ? _1541 : _1540;
    assign _1553 = ~ _1547;
    assign read_enable_70 = _102 & _1553;
    assign address_87 = _1547 ? _60 : _1529;
    assign _1549 = ~ _1547;
    assign read_enable_71 = _102 & _1549;
    assign _1547 = ~ PHASE_20;
    assign write_enable_87 = _1518 & _1547;
    assign _1551 = write_enable_87 | read_enable_71;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_42
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1551), .regcea(vdd), .wea(write_enable_87), .addra(address_87), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_70), .regceb(vdd), .web(write_enable_86), .addrb(address_86), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1558[131:131]), .sbiterrb(_1558[130:130]), .doutb(_1558[129:66]), .dbiterra(_1558[65:65]), .sbiterra(_1558[64:64]), .douta(_1558[63:0]) );
    assign _1559 = _1558[63:0];
    assign _1539 = _172[5:5];
    assign _1538 = _172[4:4];
    assign _1537 = _172[3:3];
    assign _1536 = _172[2:2];
    assign _1535 = _172[1:1];
    assign _1534 = _172[0:0];
    assign _1540 = { _1534, _1535, _1536, _1537, _1538, _1539 };
    assign address_88 = PHASE_20 ? _1541 : _1540;
    assign _1531 = ~ PHASE_20;
    assign read_enable_72 = _102 & _1531;
    assign data_85 = wr_d0;
    assign _60 = wr_addr;
    assign _1528 = _137[5:5];
    assign _1527 = _137[4:4];
    assign _1526 = _137[3:3];
    assign _1525 = _137[2:2];
    assign _1524 = _137[1:1];
    assign _1523 = _137[0:0];
    assign _1529 = { _1523, _1524, _1525, _1526, _1527, _1528 };
    assign address_89 = PHASE_20 ? _60 : _1529;
    assign _1520 = ~ PHASE_20;
    assign read_enable_73 = _102 & _1520;
    assign _62 = wr_en;
    assign _1518 = _62[0:0];
    assign write_enable_89 = _1518 & PHASE_20;
    assign _1522 = write_enable_89 | read_enable_73;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_43
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1522), .regcea(vdd), .wea(write_enable_89), .addra(address_89), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_72), .regceb(vdd), .web(write_enable_88), .addrb(address_88), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1545[131:131]), .sbiterrb(_1545[130:130]), .doutb(_1545[129:66]), .dbiterra(_1545[65:65]), .sbiterra(_1545[64:64]), .douta(_1545[63:0]) );
    assign _1546 = _1545[63:0];
    assign _1479 = ~ PHASE_20;
    assign _63 = _1479;
    always @(posedge _84) begin
        if (_82)
            PHASE_20 <= _1477;
        else
            if (_72)
                PHASE_20 <= _63;
    end
    assign _1560 = PHASE_20 ? _1559 : _1546;
    assign address_90 = _1503 ? _199 : _172;
    assign _1510 = ~ _1503;
    assign read_enable_74 = _102 & _1510;
    assign write_enable_90 = _1494 & _1503;
    assign _1512 = write_enable_90 | read_enable_74;
    assign address_91 = _1503 ? _164 : _137;
    assign _1505 = ~ _1503;
    assign read_enable_75 = _102 & _1505;
    assign _1503 = ~ PHASE_21;
    assign write_enable_91 = _1487 & _1503;
    assign _1507 = write_enable_91 | read_enable_75;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_44
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1507), .regcea(vdd), .wea(write_enable_91), .addra(address_91), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1512), .regceb(vdd), .web(write_enable_90), .addrb(address_90), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1515[131:131]), .sbiterrb(_1515[130:130]), .doutb(_1515[129:66]), .dbiterra(_1515[65:65]), .sbiterra(_1515[64:64]), .douta(_1515[63:0]) );
    assign _1516 = _1515[63:0];
    assign _1571 = _1570[127:64];
    assign data_87 = _1571;
    always @(posedge _84) begin
        if (_82)
            _175 <= _174;
        else
            _175 <= _172;
    end
    always @(posedge _84) begin
        if (_82)
            _178 <= _177;
        else
            _178 <= _175;
    end
    always @(posedge _84) begin
        if (_82)
            _181 <= _180;
        else
            _181 <= _178;
    end
    always @(posedge _84) begin
        if (_82)
            _184 <= _183;
        else
            _184 <= _181;
    end
    always @(posedge _84) begin
        if (_82)
            _187 <= _186;
        else
            _187 <= _184;
    end
    always @(posedge _84) begin
        if (_82)
            _190 <= _189;
        else
            _190 <= _187;
    end
    always @(posedge _84) begin
        if (_82)
            _193 <= _192;
        else
            _193 <= _190;
    end
    always @(posedge _84) begin
        if (_82)
            _196 <= _195;
        else
            _196 <= _193;
    end
    always @(posedge _84) begin
        if (_82)
            _199 <= _198;
        else
            _199 <= _196;
    end
    assign _172 = _91[33:28];
    assign address_92 = PHASE_21 ? _199 : _172;
    assign _1496 = ~ PHASE_21;
    assign read_enable_76 = _102 & _1496;
    assign _1493 = ~ _130;
    assign _1494 = _129 & _1493;
    assign write_enable_92 = _1494 & PHASE_21;
    assign _1498 = write_enable_92 | read_enable_76;
    assign address_93 = PHASE_21 ? _164 : _137;
    assign _1489 = ~ PHASE_21;
    assign read_enable_77 = _102 & _1489;
    assign _1486 = ~ _130;
    assign _1487 = _129 & _1486;
    assign write_enable_93 = _1487 & PHASE_21;
    assign _1491 = write_enable_93 | read_enable_77;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_45
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1491), .regcea(vdd), .wea(write_enable_93), .addra(address_93), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1498), .regceb(vdd), .web(write_enable_92), .addrb(address_92), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1501[131:131]), .sbiterrb(_1501[130:130]), .doutb(_1501[129:66]), .dbiterra(_1501[65:65]), .sbiterra(_1501[64:64]), .douta(_1501[63:0]) );
    assign _1502 = _1501[63:0];
    assign _99 = _91[492:492];
    assign _1572 = ~ PHASE_21;
    assign _65 = _1572;
    always @(posedge _84) begin
        if (_82)
            PHASE_21 <= _1484;
        else
            if (_99)
                PHASE_21 <= _65;
    end
    assign q0_6 = PHASE_21 ? _1516 : _1502;
    assign _92 = _91[483:483];
    always @(posedge _84) begin
        if (_82)
            _1482 <= _1481;
        else
            _1482 <= _92;
    end
    assign _1561 = _1482 ? _1560 : q0_6;
    dp_7
        dp
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1561), .d2(_1568), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_1570[191:128]), .q2(_1570[127:64]), .q1(_1570[63:0]) );
    assign _1573 = _1570[63:0];
    assign data_91 = _1573;
    assign _137 = _91[27:22];
    always @(posedge _84) begin
        if (_82)
            _140 <= _139;
        else
            _140 <= _137;
    end
    always @(posedge _84) begin
        if (_82)
            _143 <= _142;
        else
            _143 <= _140;
    end
    always @(posedge _84) begin
        if (_82)
            _146 <= _145;
        else
            _146 <= _143;
    end
    always @(posedge _84) begin
        if (_82)
            _149 <= _148;
        else
            _149 <= _146;
    end
    always @(posedge _84) begin
        if (_82)
            _152 <= _151;
        else
            _152 <= _149;
    end
    always @(posedge _84) begin
        if (_82)
            _155 <= _154;
        else
            _155 <= _152;
    end
    always @(posedge _84) begin
        if (_82)
            _158 <= _157;
        else
            _158 <= _155;
    end
    always @(posedge _84) begin
        if (_82)
            _161 <= _160;
        else
            _161 <= _158;
    end
    always @(posedge _84) begin
        if (_82)
            _164 <= _163;
        else
            _164 <= _161;
    end
    assign _68 = rd_addr;
    assign address_94 = PHASE_22 ? _164 : _68;
    assign _1637 = ~ PHASE_22;
    assign _70 = rd_en;
    assign _1636 = _70[0:0];
    assign read_enable_78 = _1636 & _1637;
    assign _278 = _91[485:485];
    always @(posedge _84) begin
        if (_82)
            _1607 <= _1606;
        else
            _1607 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _1610 <= _1609;
        else
            _1610 <= _1607;
    end
    always @(posedge _84) begin
        if (_82)
            _1613 <= _1612;
        else
            _1613 <= _1610;
    end
    always @(posedge _84) begin
        if (_82)
            _1616 <= _1615;
        else
            _1616 <= _1613;
    end
    always @(posedge _84) begin
        if (_82)
            _1619 <= _1618;
        else
            _1619 <= _1616;
    end
    always @(posedge _84) begin
        if (_82)
            _1622 <= _1621;
        else
            _1622 <= _1619;
    end
    always @(posedge _84) begin
        if (_82)
            _1625 <= _1624;
        else
            _1625 <= _1622;
    end
    always @(posedge _84) begin
        if (_82)
            _1628 <= _1627;
        else
            _1628 <= _1625;
    end
    always @(posedge _84) begin
        if (_82)
            _1631 <= _1630;
        else
            _1631 <= _1628;
    end
    assign _1632 = ~ _1631;
    assign _130 = _91[484:484];
    always @(posedge _84) begin
        if (_82)
            _1580 <= _1579;
        else
            _1580 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1583 <= _1582;
        else
            _1583 <= _1580;
    end
    always @(posedge _84) begin
        if (_82)
            _1586 <= _1585;
        else
            _1586 <= _1583;
    end
    always @(posedge _84) begin
        if (_82)
            _1589 <= _1588;
        else
            _1589 <= _1586;
    end
    always @(posedge _84) begin
        if (_82)
            _1592 <= _1591;
        else
            _1592 <= _1589;
    end
    always @(posedge _84) begin
        if (_82)
            _1595 <= _1594;
        else
            _1595 <= _1592;
    end
    always @(posedge _84) begin
        if (_82)
            _1598 <= _1597;
        else
            _1598 <= _1595;
    end
    always @(posedge _84) begin
        if (_82)
            _1601 <= _1600;
        else
            _1601 <= _1598;
    end
    always @(posedge _84) begin
        if (_82)
            _1604 <= _1603;
        else
            _1604 <= _1601;
    end
    assign _1633 = _1604 & _1632;
    assign _102 = _91[491:491];
    always @(posedge _84) begin
        if (_82)
            _105 <= _104;
        else
            _105 <= _102;
    end
    always @(posedge _84) begin
        if (_82)
            _108 <= _107;
        else
            _108 <= _105;
    end
    always @(posedge _84) begin
        if (_82)
            _111 <= _110;
        else
            _111 <= _108;
    end
    always @(posedge _84) begin
        if (_82)
            _114 <= _113;
        else
            _114 <= _111;
    end
    always @(posedge _84) begin
        if (_82)
            _117 <= _116;
        else
            _117 <= _114;
    end
    always @(posedge _84) begin
        if (_82)
            _120 <= _119;
        else
            _120 <= _117;
    end
    always @(posedge _84) begin
        if (_82)
            _123 <= _122;
        else
            _123 <= _120;
    end
    always @(posedge _84) begin
        if (_82)
            _126 <= _125;
        else
            _126 <= _123;
    end
    always @(posedge _84) begin
        if (_82)
            _129 <= _128;
        else
            _129 <= _126;
    end
    assign _1634 = _129 & _1633;
    assign write_enable_94 = _1634 & PHASE_22;
    assign _1639 = write_enable_94 | read_enable_78;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_46
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1639), .regcea(vdd), .wea(write_enable_94), .addra(address_94), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_85), .regceb(vdd), .web(write_enable_85), .addrb(address_85), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1646[131:131]), .sbiterrb(_1646[130:130]), .doutb(_1646[129:66]), .dbiterra(_1646[65:65]), .sbiterra(_1646[64:64]), .douta(_1646[63:0]) );
    assign _1647 = _1646[63:0];
    assign _72 = flip;
    assign _1577 = ~ PHASE_22;
    assign _73 = _1577;
    always @(posedge _84) begin
        if (_82)
            PHASE_22 <= _1575;
        else
            if (_72)
                PHASE_22 <= _73;
    end
    assign _1659 = PHASE_22 ? _1658 : _1647;
    assign _76 = first_4step_pass;
    assign _78 = first_iter;
    assign _80 = start;
    assign _82 = clear;
    assign _84 = clock;
    ctrl
        ctrl
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .first_4step_pass(_76), .flip(_91[492:492]), .read_write_enable(_91[491:491]), .index(_91[490:487]), .valid(_91[486:486]), .twiddle_stage(_91[485:485]), .last_stage(_91[484:484]), .first_stage(_91[483:483]), .start_twiddles(_91[482:482]), .omegas6(_91[481:418]), .omegas5(_91[417:354]), .omegas4(_91[353:290]), .omegas3(_91[289:226]), .omegas2(_91[225:162]), .omegas1(_91[161:98]), .omegas0(_91[97:34]), .addr2(_91[33:28]), .addr1(_91[27:22]), .m(_91[21:16]), .k(_91[15:10]), .j(_91[9:4]), .i(_91[3:1]), .done_(_91[0:0]) );
    assign _1660 = _91[0:0];

    /* aliases */
    assign data_0 = data;
    assign data_2 = data_1;
    assign data_4 = data_3;
    assign data_5 = data_3;
    assign data_6 = data_3;
    assign data_8 = data_7;
    assign data_9 = data_7;
    assign data_10 = data_7;
    assign data_12 = data_11;
    assign data_14 = data_13;
    assign data_16 = data_15;
    assign data_17 = data_15;
    assign data_18 = data_15;
    assign data_20 = data_19;
    assign data_21 = data_19;
    assign data_22 = data_19;
    assign data_24 = data_23;
    assign data_26 = data_25;
    assign data_28 = data_27;
    assign data_29 = data_27;
    assign data_30 = data_27;
    assign data_32 = data_31;
    assign data_33 = data_31;
    assign data_34 = data_31;
    assign data_36 = data_35;
    assign data_38 = data_37;
    assign data_40 = data_39;
    assign data_41 = data_39;
    assign data_42 = data_39;
    assign data_44 = data_43;
    assign data_45 = data_43;
    assign data_46 = data_43;
    assign data_48 = data_47;
    assign data_50 = data_49;
    assign data_52 = data_51;
    assign data_53 = data_51;
    assign data_54 = data_51;
    assign data_56 = data_55;
    assign data_57 = data_55;
    assign data_58 = data_55;
    assign data_60 = data_59;
    assign data_62 = data_61;
    assign data_64 = data_63;
    assign data_65 = data_63;
    assign data_66 = data_63;
    assign data_68 = data_67;
    assign data_69 = data_67;
    assign data_70 = data_67;
    assign data_72 = data_71;
    assign data_74 = data_73;
    assign data_76 = data_75;
    assign data_77 = data_75;
    assign data_78 = data_75;
    assign data_80 = data_79;
    assign data_81 = data_79;
    assign data_82 = data_79;
    assign data_84 = data_83;
    assign data_86 = data_85;
    assign data_88 = data_87;
    assign data_89 = data_87;
    assign data_90 = data_87;
    assign data_92 = data_91;
    assign data_93 = data_91;
    assign data_94 = data_91;

    /* output assignments */
    assign done_ = _1660;
    assign rd_q0 = _1659;
    assign rd_q1 = _1475;
    assign rd_q2 = _1291;
    assign rd_q3 = _1107;
    assign rd_q4 = _923;
    assign rd_q5 = _739;
    assign rd_q6 = _555;
    assign rd_q7 = _371;

endmodule
module dp_15 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0011101110101011111110001010011100001011100100000001011011010111;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1100001011011110110100010111001001000011011101011110000100101110;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0000001111101000110111111101001001001110100011100111100000011111;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1011111101111001000101000011110011100110000011001010100101100110;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_16 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1111101001000001000010100110000110101001010000001100100110010001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0011101110111001101010001100100111100110111001100010110110000001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0000101011010100001111101101111100000110100100101100100100101100;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1100011100000010001001001100010100111000011010101001001111101100;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1000010101101100110100111011111111110010000000100110100111010001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0011010000011101000101101001000011011011010010010000110100100111;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0100100110100010100000100001010001100101001101010001011100011101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_17 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0011100101000011001000100101011011000011001110101010011001010110;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1010100110001010110101010011000100100110101001101111101110101001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0111001100001110001111011101000101111010000101110111100100101011;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1010001101110111101111000010110101111101000101111110101011000110;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0111010010100011111001001101111110000010101010011101010011011100;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1110010100001110110001011011010111010011000010010011010110000000;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0011101010100111000001000000100000001000111011011010110011010101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_18 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0001010111001101000110011110110000111000111011000110110011000000;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1100000110100101110110001101011101010001111011111100110000101001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1010010100110011110001111100101101100000101100110000011111111100;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1000101100001010111010001010110010111101100011001011110110100011;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1000001111111001000110011011011001110010101010001001011001000010;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0110101000110010001100111010010010010100010001010011111110101101;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0111110110111110000110111110000001011100001011100001001111111100;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_19 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0100101111010011001001111101111001111010100010111010100101011100;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0101101010011100111100001000011100111110010010010000110000101110;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0000101111111101100110101110100101111000100111010010010010100100;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1100001011011110110100010111001001000011011101011110000100101110;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0011100110101111101011010110110000110010100010110001011011110110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1100100001000011111100010110001010010100011000001011010101010001;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0011110110100000010111111110111001110000110001001111001010111010;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_20 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1000010011111110111000001000111111110100000010001110100011110101;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0011100101000011001000100101011011000011001110101010011001010110;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0100110101000101100110100100101010000010100001001110100110001011;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0011001010101001010101000011100000101111110100000000100010101001;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0101011011000110011100011000111110000111111100001101111000100011;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0110110110111110101101111110000000100110100001110010111000111001;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1110100111110010110110100110110010111110001000101100111000010001;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_21 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1001001011011011011111100011110001111000111000010001011100001010;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1011011001011100010110001001101101111110111011011001110100000001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0011101000011111001001000011010101011110111100010101101111011100;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1101111001111011001000111110011111101101000010100101000100111011;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1111101010111110101001111000110111010110001001011011111111101111;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0100101110110010101100100000100001100011101000000110001110100010;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1010111010000110001000110110000101111000100111001100001010010101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_22 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0000011011101000101001110111110111010011010010001110011101111000;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0000100111111001111000010110100110110000101000001000011001100001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1011011110011110110010000111100001001001100101100001111111000101;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0010011111110000100011101111111110010100001010001111010101010110;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1010011110001110001001110010010111011000100111010111001100001110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1101110101000010000111010100011101101011001100100010000100000001;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1000100110001011100100100101110100111011001111100011100111000111;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module parallel_cores_1 (
    wr_d7,
    wr_d6,
    wr_d5,
    wr_d4,
    wr_d3,
    wr_d2,
    wr_d1,
    wr_d0,
    wr_addr,
    wr_en,
    rd_addr,
    rd_en,
    flip,
    first_4step_pass,
    first_iter,
    start,
    clear,
    clock,
    done_,
    rd_q0,
    rd_q1,
    rd_q2,
    rd_q3,
    rd_q4,
    rd_q5,
    rd_q6,
    rd_q7
);

    input [63:0] wr_d7;
    input [63:0] wr_d6;
    input [63:0] wr_d5;
    input [63:0] wr_d4;
    input [63:0] wr_d3;
    input [63:0] wr_d2;
    input [63:0] wr_d1;
    input [63:0] wr_d0;
    input [5:0] wr_addr;
    input [7:0] wr_en;
    input [5:0] rd_addr;
    input [7:0] rd_en;
    input flip;
    input first_4step_pass;
    input first_iter;
    input start;
    input clear;
    input clock;
    output done_;
    output [63:0] rd_q0;
    output [63:0] rd_q1;
    output [63:0] rd_q2;
    output [63:0] rd_q3;
    output [63:0] rd_q4;
    output [63:0] rd_q5;
    output [63:0] rd_q6;
    output [63:0] rd_q7;

    /* signal declarations */
    wire [5:0] address;
    wire write_enable;
    wire [5:0] address_0;
    wire _362;
    wire read_enable;
    wire _360;
    wire write_enable_0;
    wire _364;
    wire [131:0] _369;
    wire [63:0] _370;
    wire [5:0] _355 = 6'b000000;
    wire [5:0] address_1;
    wire _353;
    wire write_enable_1;
    wire [63:0] _267;
    wire [63:0] _266;
    wire [63:0] _268;
    wire [63:0] _264;
    wire [63:0] _263;
    wire [63:0] q1;
    wire [63:0] _269;
    wire [5:0] address_2;
    wire write_enable_2 = 1'b0;
    wire _254;
    wire read_enable_0;
    wire [5:0] address_3;
    wire _250;
    wire read_enable_1;
    wire _248;
    wire write_enable_3;
    wire _252;
    wire [131:0] _259;
    wire [63:0] _260;
    wire [63:0] data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_0;
    wire [5:0] _242 = 6'b000000;
    wire _240;
    wire _239;
    wire _238;
    wire _237;
    wire _236;
    wire _235;
    wire [5:0] _241;
    wire [5:0] address_4;
    wire write_enable_4 = 1'b0;
    wire _232;
    wire read_enable_2;
    wire [63:0] data_1;
    wire [63:0] data_2;
    wire _229;
    wire _228;
    wire _227;
    wire _226;
    wire _225;
    wire _224;
    wire [5:0] _230;
    wire [5:0] address_5;
    wire _221;
    wire read_enable_3;
    wire _219;
    wire write_enable_5;
    wire _223;
    wire [131:0] _246;
    wire [63:0] _247;
    wire _87 = 1'b0;
    wire _86 = 1'b0;
    wire _89;
    wire _3;
    reg PHASE;
    wire [63:0] _261;
    wire [5:0] address_6;
    wire _211;
    wire read_enable_4;
    wire write_enable_6;
    wire _213;
    wire [5:0] address_7;
    wire _206;
    wire read_enable_5;
    wire _204;
    wire write_enable_7;
    wire _208;
    wire [131:0] _216;
    wire [63:0] _217;
    wire [63:0] _283;
    wire [63:0] data_3;
    wire [63:0] data_4;
    wire [63:0] data_5;
    wire [63:0] data_6;
    wire [5:0] address_8;
    wire _169;
    wire read_enable_6;
    wire _166;
    wire _167;
    wire write_enable_8;
    wire _171;
    wire [5:0] address_9;
    wire _134;
    wire read_enable_7;
    wire _131;
    wire _132;
    wire write_enable_9;
    wire _136;
    wire [131:0] _202;
    wire [63:0] _203;
    wire _98 = 1'b0;
    wire _97 = 1'b0;
    wire _284;
    wire _5;
    reg PHASE_0;
    wire [63:0] q0;
    wire _94 = 1'b0;
    wire _93 = 1'b0;
    reg _96;
    wire [63:0] _262;
    wire [191:0] _282;
    wire [63:0] _285;
    wire [63:0] data_7;
    wire [63:0] data_8;
    wire [63:0] data_9;
    wire [63:0] data_10;
    wire [5:0] address_10;
    wire _349;
    wire _348;
    wire read_enable_8;
    wire _342 = 1'b0;
    wire _341 = 1'b0;
    wire _339 = 1'b0;
    wire _338 = 1'b0;
    wire _336 = 1'b0;
    wire _335 = 1'b0;
    wire _333 = 1'b0;
    wire _332 = 1'b0;
    wire _330 = 1'b0;
    wire _329 = 1'b0;
    wire _327 = 1'b0;
    wire _326 = 1'b0;
    wire _324 = 1'b0;
    wire _323 = 1'b0;
    wire _321 = 1'b0;
    wire _320 = 1'b0;
    wire _318 = 1'b0;
    wire _317 = 1'b0;
    reg _319;
    reg _322;
    reg _325;
    reg _328;
    reg _331;
    reg _334;
    reg _337;
    reg _340;
    reg _343;
    wire _344;
    wire _315 = 1'b0;
    wire _314 = 1'b0;
    wire _312 = 1'b0;
    wire _311 = 1'b0;
    wire _309 = 1'b0;
    wire _308 = 1'b0;
    wire _306 = 1'b0;
    wire _305 = 1'b0;
    wire _303 = 1'b0;
    wire _302 = 1'b0;
    wire _300 = 1'b0;
    wire _299 = 1'b0;
    wire _297 = 1'b0;
    wire _296 = 1'b0;
    wire _294 = 1'b0;
    wire _293 = 1'b0;
    wire _291 = 1'b0;
    wire _290 = 1'b0;
    reg _292;
    reg _295;
    reg _298;
    reg _301;
    reg _304;
    reg _307;
    reg _310;
    reg _313;
    reg _316;
    wire _345;
    wire _346;
    wire write_enable_10;
    wire _351;
    wire [131:0] _358;
    wire [63:0] _359;
    wire _287 = 1'b0;
    wire _286 = 1'b0;
    wire _289;
    wire _7;
    reg PHASE_1;
    wire [63:0] _371;
    wire [5:0] address_11;
    wire write_enable_11;
    wire [5:0] address_12;
    wire _546;
    wire read_enable_9;
    wire _544;
    wire write_enable_12;
    wire _548;
    wire [131:0] _553;
    wire [63:0] _554;
    wire [5:0] _539 = 6'b000000;
    wire [5:0] address_13;
    wire _537;
    wire write_enable_13;
    wire [63:0] _462;
    wire [63:0] _461;
    wire [63:0] _463;
    wire [63:0] _459;
    wire [63:0] _458;
    wire [63:0] q1_0;
    wire [63:0] _464;
    wire [5:0] address_14;
    wire write_enable_14 = 1'b0;
    wire _449;
    wire read_enable_10;
    wire [5:0] address_15;
    wire _445;
    wire read_enable_11;
    wire _443;
    wire write_enable_15;
    wire _447;
    wire [131:0] _454;
    wire [63:0] _455;
    wire [63:0] data_11 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_12;
    wire [5:0] _437 = 6'b000000;
    wire _435;
    wire _434;
    wire _433;
    wire _432;
    wire _431;
    wire _430;
    wire [5:0] _436;
    wire [5:0] address_16;
    wire write_enable_16 = 1'b0;
    wire _427;
    wire read_enable_12;
    wire [63:0] data_13;
    wire [63:0] data_14;
    wire _424;
    wire _423;
    wire _422;
    wire _421;
    wire _420;
    wire _419;
    wire [5:0] _425;
    wire [5:0] address_17;
    wire _416;
    wire read_enable_13;
    wire _414;
    wire write_enable_17;
    wire _418;
    wire [131:0] _441;
    wire [63:0] _442;
    wire _373 = 1'b0;
    wire _372 = 1'b0;
    wire _375;
    wire _11;
    reg PHASE_2;
    wire [63:0] _456;
    wire [5:0] address_18;
    wire _406;
    wire read_enable_14;
    wire write_enable_18;
    wire _408;
    wire [5:0] address_19;
    wire _401;
    wire read_enable_15;
    wire _399;
    wire write_enable_19;
    wire _403;
    wire [131:0] _411;
    wire [63:0] _412;
    wire [63:0] _467;
    wire [63:0] data_15;
    wire [63:0] data_16;
    wire [63:0] data_17;
    wire [63:0] data_18;
    wire [5:0] address_20;
    wire _392;
    wire read_enable_16;
    wire _389;
    wire _390;
    wire write_enable_20;
    wire _394;
    wire [5:0] address_21;
    wire _385;
    wire read_enable_17;
    wire _382;
    wire _383;
    wire write_enable_21;
    wire _387;
    wire [131:0] _397;
    wire [63:0] _398;
    wire _380 = 1'b0;
    wire _379 = 1'b0;
    wire _468;
    wire _13;
    reg PHASE_3;
    wire [63:0] q0_0;
    wire _377 = 1'b0;
    wire _376 = 1'b0;
    reg _378;
    wire [63:0] _457;
    wire [191:0] _466;
    wire [63:0] _469;
    wire [63:0] data_19;
    wire [63:0] data_20;
    wire [63:0] data_21;
    wire [63:0] data_22;
    wire [5:0] address_22;
    wire _533;
    wire _532;
    wire read_enable_18;
    wire _526 = 1'b0;
    wire _525 = 1'b0;
    wire _523 = 1'b0;
    wire _522 = 1'b0;
    wire _520 = 1'b0;
    wire _519 = 1'b0;
    wire _517 = 1'b0;
    wire _516 = 1'b0;
    wire _514 = 1'b0;
    wire _513 = 1'b0;
    wire _511 = 1'b0;
    wire _510 = 1'b0;
    wire _508 = 1'b0;
    wire _507 = 1'b0;
    wire _505 = 1'b0;
    wire _504 = 1'b0;
    wire _502 = 1'b0;
    wire _501 = 1'b0;
    reg _503;
    reg _506;
    reg _509;
    reg _512;
    reg _515;
    reg _518;
    reg _521;
    reg _524;
    reg _527;
    wire _528;
    wire _499 = 1'b0;
    wire _498 = 1'b0;
    wire _496 = 1'b0;
    wire _495 = 1'b0;
    wire _493 = 1'b0;
    wire _492 = 1'b0;
    wire _490 = 1'b0;
    wire _489 = 1'b0;
    wire _487 = 1'b0;
    wire _486 = 1'b0;
    wire _484 = 1'b0;
    wire _483 = 1'b0;
    wire _481 = 1'b0;
    wire _480 = 1'b0;
    wire _478 = 1'b0;
    wire _477 = 1'b0;
    wire _475 = 1'b0;
    wire _474 = 1'b0;
    reg _476;
    reg _479;
    reg _482;
    reg _485;
    reg _488;
    reg _491;
    reg _494;
    reg _497;
    reg _500;
    wire _529;
    wire _530;
    wire write_enable_22;
    wire _535;
    wire [131:0] _542;
    wire [63:0] _543;
    wire _471 = 1'b0;
    wire _470 = 1'b0;
    wire _473;
    wire _15;
    reg PHASE_4;
    wire [63:0] _555;
    wire [5:0] address_23;
    wire write_enable_23;
    wire [5:0] address_24;
    wire _730;
    wire read_enable_19;
    wire _728;
    wire write_enable_24;
    wire _732;
    wire [131:0] _737;
    wire [63:0] _738;
    wire [5:0] _723 = 6'b000000;
    wire [5:0] address_25;
    wire _721;
    wire write_enable_25;
    wire [63:0] _646;
    wire [63:0] _645;
    wire [63:0] _647;
    wire [63:0] _643;
    wire [63:0] _642;
    wire [63:0] q1_1;
    wire [63:0] _648;
    wire [5:0] address_26;
    wire write_enable_26 = 1'b0;
    wire _633;
    wire read_enable_20;
    wire [5:0] address_27;
    wire _629;
    wire read_enable_21;
    wire _627;
    wire write_enable_27;
    wire _631;
    wire [131:0] _638;
    wire [63:0] _639;
    wire [63:0] data_23 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_24;
    wire [5:0] _621 = 6'b000000;
    wire _619;
    wire _618;
    wire _617;
    wire _616;
    wire _615;
    wire _614;
    wire [5:0] _620;
    wire [5:0] address_28;
    wire write_enable_28 = 1'b0;
    wire _611;
    wire read_enable_22;
    wire [63:0] data_25;
    wire [63:0] data_26;
    wire _608;
    wire _607;
    wire _606;
    wire _605;
    wire _604;
    wire _603;
    wire [5:0] _609;
    wire [5:0] address_29;
    wire _600;
    wire read_enable_23;
    wire _598;
    wire write_enable_29;
    wire _602;
    wire [131:0] _625;
    wire [63:0] _626;
    wire _557 = 1'b0;
    wire _556 = 1'b0;
    wire _559;
    wire _19;
    reg PHASE_5;
    wire [63:0] _640;
    wire [5:0] address_30;
    wire _590;
    wire read_enable_24;
    wire write_enable_30;
    wire _592;
    wire [5:0] address_31;
    wire _585;
    wire read_enable_25;
    wire _583;
    wire write_enable_31;
    wire _587;
    wire [131:0] _595;
    wire [63:0] _596;
    wire [63:0] _651;
    wire [63:0] data_27;
    wire [63:0] data_28;
    wire [63:0] data_29;
    wire [63:0] data_30;
    wire [5:0] address_32;
    wire _576;
    wire read_enable_26;
    wire _573;
    wire _574;
    wire write_enable_32;
    wire _578;
    wire [5:0] address_33;
    wire _569;
    wire read_enable_27;
    wire _566;
    wire _567;
    wire write_enable_33;
    wire _571;
    wire [131:0] _581;
    wire [63:0] _582;
    wire _564 = 1'b0;
    wire _563 = 1'b0;
    wire _652;
    wire _21;
    reg PHASE_6;
    wire [63:0] q0_1;
    wire _561 = 1'b0;
    wire _560 = 1'b0;
    reg _562;
    wire [63:0] _641;
    wire [191:0] _650;
    wire [63:0] _653;
    wire [63:0] data_31;
    wire [63:0] data_32;
    wire [63:0] data_33;
    wire [63:0] data_34;
    wire [5:0] address_34;
    wire _717;
    wire _716;
    wire read_enable_28;
    wire _710 = 1'b0;
    wire _709 = 1'b0;
    wire _707 = 1'b0;
    wire _706 = 1'b0;
    wire _704 = 1'b0;
    wire _703 = 1'b0;
    wire _701 = 1'b0;
    wire _700 = 1'b0;
    wire _698 = 1'b0;
    wire _697 = 1'b0;
    wire _695 = 1'b0;
    wire _694 = 1'b0;
    wire _692 = 1'b0;
    wire _691 = 1'b0;
    wire _689 = 1'b0;
    wire _688 = 1'b0;
    wire _686 = 1'b0;
    wire _685 = 1'b0;
    reg _687;
    reg _690;
    reg _693;
    reg _696;
    reg _699;
    reg _702;
    reg _705;
    reg _708;
    reg _711;
    wire _712;
    wire _683 = 1'b0;
    wire _682 = 1'b0;
    wire _680 = 1'b0;
    wire _679 = 1'b0;
    wire _677 = 1'b0;
    wire _676 = 1'b0;
    wire _674 = 1'b0;
    wire _673 = 1'b0;
    wire _671 = 1'b0;
    wire _670 = 1'b0;
    wire _668 = 1'b0;
    wire _667 = 1'b0;
    wire _665 = 1'b0;
    wire _664 = 1'b0;
    wire _662 = 1'b0;
    wire _661 = 1'b0;
    wire _659 = 1'b0;
    wire _658 = 1'b0;
    reg _660;
    reg _663;
    reg _666;
    reg _669;
    reg _672;
    reg _675;
    reg _678;
    reg _681;
    reg _684;
    wire _713;
    wire _714;
    wire write_enable_34;
    wire _719;
    wire [131:0] _726;
    wire [63:0] _727;
    wire _655 = 1'b0;
    wire _654 = 1'b0;
    wire _657;
    wire _23;
    reg PHASE_7;
    wire [63:0] _739;
    wire [5:0] address_35;
    wire write_enable_35;
    wire [5:0] address_36;
    wire _914;
    wire read_enable_29;
    wire _912;
    wire write_enable_36;
    wire _916;
    wire [131:0] _921;
    wire [63:0] _922;
    wire [5:0] _907 = 6'b000000;
    wire [5:0] address_37;
    wire _905;
    wire write_enable_37;
    wire [63:0] _830;
    wire [63:0] _829;
    wire [63:0] _831;
    wire [63:0] _827;
    wire [63:0] _826;
    wire [63:0] q1_2;
    wire [63:0] _832;
    wire [5:0] address_38;
    wire write_enable_38 = 1'b0;
    wire _817;
    wire read_enable_30;
    wire [5:0] address_39;
    wire _813;
    wire read_enable_31;
    wire _811;
    wire write_enable_39;
    wire _815;
    wire [131:0] _822;
    wire [63:0] _823;
    wire [63:0] data_35 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_36;
    wire [5:0] _805 = 6'b000000;
    wire _803;
    wire _802;
    wire _801;
    wire _800;
    wire _799;
    wire _798;
    wire [5:0] _804;
    wire [5:0] address_40;
    wire write_enable_40 = 1'b0;
    wire _795;
    wire read_enable_32;
    wire [63:0] data_37;
    wire [63:0] data_38;
    wire _792;
    wire _791;
    wire _790;
    wire _789;
    wire _788;
    wire _787;
    wire [5:0] _793;
    wire [5:0] address_41;
    wire _784;
    wire read_enable_33;
    wire _782;
    wire write_enable_41;
    wire _786;
    wire [131:0] _809;
    wire [63:0] _810;
    wire _741 = 1'b0;
    wire _740 = 1'b0;
    wire _743;
    wire _27;
    reg PHASE_8;
    wire [63:0] _824;
    wire [5:0] address_42;
    wire _774;
    wire read_enable_34;
    wire write_enable_42;
    wire _776;
    wire [5:0] address_43;
    wire _769;
    wire read_enable_35;
    wire _767;
    wire write_enable_43;
    wire _771;
    wire [131:0] _779;
    wire [63:0] _780;
    wire [63:0] _835;
    wire [63:0] data_39;
    wire [63:0] data_40;
    wire [63:0] data_41;
    wire [63:0] data_42;
    wire [5:0] address_44;
    wire _760;
    wire read_enable_36;
    wire _757;
    wire _758;
    wire write_enable_44;
    wire _762;
    wire [5:0] address_45;
    wire _753;
    wire read_enable_37;
    wire _750;
    wire _751;
    wire write_enable_45;
    wire _755;
    wire [131:0] _765;
    wire [63:0] _766;
    wire _748 = 1'b0;
    wire _747 = 1'b0;
    wire _836;
    wire _29;
    reg PHASE_9;
    wire [63:0] q0_2;
    wire _745 = 1'b0;
    wire _744 = 1'b0;
    reg _746;
    wire [63:0] _825;
    wire [191:0] _834;
    wire [63:0] _837;
    wire [63:0] data_43;
    wire [63:0] data_44;
    wire [63:0] data_45;
    wire [63:0] data_46;
    wire [5:0] address_46;
    wire _901;
    wire _900;
    wire read_enable_38;
    wire _894 = 1'b0;
    wire _893 = 1'b0;
    wire _891 = 1'b0;
    wire _890 = 1'b0;
    wire _888 = 1'b0;
    wire _887 = 1'b0;
    wire _885 = 1'b0;
    wire _884 = 1'b0;
    wire _882 = 1'b0;
    wire _881 = 1'b0;
    wire _879 = 1'b0;
    wire _878 = 1'b0;
    wire _876 = 1'b0;
    wire _875 = 1'b0;
    wire _873 = 1'b0;
    wire _872 = 1'b0;
    wire _870 = 1'b0;
    wire _869 = 1'b0;
    reg _871;
    reg _874;
    reg _877;
    reg _880;
    reg _883;
    reg _886;
    reg _889;
    reg _892;
    reg _895;
    wire _896;
    wire _867 = 1'b0;
    wire _866 = 1'b0;
    wire _864 = 1'b0;
    wire _863 = 1'b0;
    wire _861 = 1'b0;
    wire _860 = 1'b0;
    wire _858 = 1'b0;
    wire _857 = 1'b0;
    wire _855 = 1'b0;
    wire _854 = 1'b0;
    wire _852 = 1'b0;
    wire _851 = 1'b0;
    wire _849 = 1'b0;
    wire _848 = 1'b0;
    wire _846 = 1'b0;
    wire _845 = 1'b0;
    wire _843 = 1'b0;
    wire _842 = 1'b0;
    reg _844;
    reg _847;
    reg _850;
    reg _853;
    reg _856;
    reg _859;
    reg _862;
    reg _865;
    reg _868;
    wire _897;
    wire _898;
    wire write_enable_46;
    wire _903;
    wire [131:0] _910;
    wire [63:0] _911;
    wire _839 = 1'b0;
    wire _838 = 1'b0;
    wire _841;
    wire _31;
    reg PHASE_10;
    wire [63:0] _923;
    wire [5:0] address_47;
    wire write_enable_47;
    wire [5:0] address_48;
    wire _1098;
    wire read_enable_39;
    wire _1096;
    wire write_enable_48;
    wire _1100;
    wire [131:0] _1105;
    wire [63:0] _1106;
    wire [5:0] _1091 = 6'b000000;
    wire [5:0] address_49;
    wire _1089;
    wire write_enable_49;
    wire [63:0] _1014;
    wire [63:0] _1013;
    wire [63:0] _1015;
    wire [63:0] _1011;
    wire [63:0] _1010;
    wire [63:0] q1_3;
    wire [63:0] _1016;
    wire [5:0] address_50;
    wire write_enable_50 = 1'b0;
    wire _1001;
    wire read_enable_40;
    wire [5:0] address_51;
    wire _997;
    wire read_enable_41;
    wire _995;
    wire write_enable_51;
    wire _999;
    wire [131:0] _1006;
    wire [63:0] _1007;
    wire [63:0] data_47 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_48;
    wire [5:0] _989 = 6'b000000;
    wire _987;
    wire _986;
    wire _985;
    wire _984;
    wire _983;
    wire _982;
    wire [5:0] _988;
    wire [5:0] address_52;
    wire write_enable_52 = 1'b0;
    wire _979;
    wire read_enable_42;
    wire [63:0] data_49;
    wire [63:0] data_50;
    wire _976;
    wire _975;
    wire _974;
    wire _973;
    wire _972;
    wire _971;
    wire [5:0] _977;
    wire [5:0] address_53;
    wire _968;
    wire read_enable_43;
    wire _966;
    wire write_enable_53;
    wire _970;
    wire [131:0] _993;
    wire [63:0] _994;
    wire _925 = 1'b0;
    wire _924 = 1'b0;
    wire _927;
    wire _35;
    reg PHASE_11;
    wire [63:0] _1008;
    wire [5:0] address_54;
    wire _958;
    wire read_enable_44;
    wire write_enable_54;
    wire _960;
    wire [5:0] address_55;
    wire _953;
    wire read_enable_45;
    wire _951;
    wire write_enable_55;
    wire _955;
    wire [131:0] _963;
    wire [63:0] _964;
    wire [63:0] _1019;
    wire [63:0] data_51;
    wire [63:0] data_52;
    wire [63:0] data_53;
    wire [63:0] data_54;
    wire [5:0] address_56;
    wire _944;
    wire read_enable_46;
    wire _941;
    wire _942;
    wire write_enable_56;
    wire _946;
    wire [5:0] address_57;
    wire _937;
    wire read_enable_47;
    wire _934;
    wire _935;
    wire write_enable_57;
    wire _939;
    wire [131:0] _949;
    wire [63:0] _950;
    wire _932 = 1'b0;
    wire _931 = 1'b0;
    wire _1020;
    wire _37;
    reg PHASE_12;
    wire [63:0] q0_3;
    wire _929 = 1'b0;
    wire _928 = 1'b0;
    reg _930;
    wire [63:0] _1009;
    wire [191:0] _1018;
    wire [63:0] _1021;
    wire [63:0] data_55;
    wire [63:0] data_56;
    wire [63:0] data_57;
    wire [63:0] data_58;
    wire [5:0] address_58;
    wire _1085;
    wire _1084;
    wire read_enable_48;
    wire _1078 = 1'b0;
    wire _1077 = 1'b0;
    wire _1075 = 1'b0;
    wire _1074 = 1'b0;
    wire _1072 = 1'b0;
    wire _1071 = 1'b0;
    wire _1069 = 1'b0;
    wire _1068 = 1'b0;
    wire _1066 = 1'b0;
    wire _1065 = 1'b0;
    wire _1063 = 1'b0;
    wire _1062 = 1'b0;
    wire _1060 = 1'b0;
    wire _1059 = 1'b0;
    wire _1057 = 1'b0;
    wire _1056 = 1'b0;
    wire _1054 = 1'b0;
    wire _1053 = 1'b0;
    reg _1055;
    reg _1058;
    reg _1061;
    reg _1064;
    reg _1067;
    reg _1070;
    reg _1073;
    reg _1076;
    reg _1079;
    wire _1080;
    wire _1051 = 1'b0;
    wire _1050 = 1'b0;
    wire _1048 = 1'b0;
    wire _1047 = 1'b0;
    wire _1045 = 1'b0;
    wire _1044 = 1'b0;
    wire _1042 = 1'b0;
    wire _1041 = 1'b0;
    wire _1039 = 1'b0;
    wire _1038 = 1'b0;
    wire _1036 = 1'b0;
    wire _1035 = 1'b0;
    wire _1033 = 1'b0;
    wire _1032 = 1'b0;
    wire _1030 = 1'b0;
    wire _1029 = 1'b0;
    wire _1027 = 1'b0;
    wire _1026 = 1'b0;
    reg _1028;
    reg _1031;
    reg _1034;
    reg _1037;
    reg _1040;
    reg _1043;
    reg _1046;
    reg _1049;
    reg _1052;
    wire _1081;
    wire _1082;
    wire write_enable_58;
    wire _1087;
    wire [131:0] _1094;
    wire [63:0] _1095;
    wire _1023 = 1'b0;
    wire _1022 = 1'b0;
    wire _1025;
    wire _39;
    reg PHASE_13;
    wire [63:0] _1107;
    wire [5:0] address_59;
    wire write_enable_59;
    wire [5:0] address_60;
    wire _1282;
    wire read_enable_49;
    wire _1280;
    wire write_enable_60;
    wire _1284;
    wire [131:0] _1289;
    wire [63:0] _1290;
    wire [5:0] _1275 = 6'b000000;
    wire [5:0] address_61;
    wire _1273;
    wire write_enable_61;
    wire [63:0] _1198;
    wire [63:0] _1197;
    wire [63:0] _1199;
    wire [63:0] _1195;
    wire [63:0] _1194;
    wire [63:0] q1_4;
    wire [63:0] _1200;
    wire [5:0] address_62;
    wire write_enable_62 = 1'b0;
    wire _1185;
    wire read_enable_50;
    wire [5:0] address_63;
    wire _1181;
    wire read_enable_51;
    wire _1179;
    wire write_enable_63;
    wire _1183;
    wire [131:0] _1190;
    wire [63:0] _1191;
    wire [63:0] data_59 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_60;
    wire [5:0] _1173 = 6'b000000;
    wire _1171;
    wire _1170;
    wire _1169;
    wire _1168;
    wire _1167;
    wire _1166;
    wire [5:0] _1172;
    wire [5:0] address_64;
    wire write_enable_64 = 1'b0;
    wire _1163;
    wire read_enable_52;
    wire [63:0] data_61;
    wire [63:0] data_62;
    wire _1160;
    wire _1159;
    wire _1158;
    wire _1157;
    wire _1156;
    wire _1155;
    wire [5:0] _1161;
    wire [5:0] address_65;
    wire _1152;
    wire read_enable_53;
    wire _1150;
    wire write_enable_65;
    wire _1154;
    wire [131:0] _1177;
    wire [63:0] _1178;
    wire _1109 = 1'b0;
    wire _1108 = 1'b0;
    wire _1111;
    wire _43;
    reg PHASE_14;
    wire [63:0] _1192;
    wire [5:0] address_66;
    wire _1142;
    wire read_enable_54;
    wire write_enable_66;
    wire _1144;
    wire [5:0] address_67;
    wire _1137;
    wire read_enable_55;
    wire _1135;
    wire write_enable_67;
    wire _1139;
    wire [131:0] _1147;
    wire [63:0] _1148;
    wire [63:0] _1203;
    wire [63:0] data_63;
    wire [63:0] data_64;
    wire [63:0] data_65;
    wire [63:0] data_66;
    wire [5:0] address_68;
    wire _1128;
    wire read_enable_56;
    wire _1125;
    wire _1126;
    wire write_enable_68;
    wire _1130;
    wire [5:0] address_69;
    wire _1121;
    wire read_enable_57;
    wire _1118;
    wire _1119;
    wire write_enable_69;
    wire _1123;
    wire [131:0] _1133;
    wire [63:0] _1134;
    wire _1116 = 1'b0;
    wire _1115 = 1'b0;
    wire _1204;
    wire _45;
    reg PHASE_15;
    wire [63:0] q0_4;
    wire _1113 = 1'b0;
    wire _1112 = 1'b0;
    reg _1114;
    wire [63:0] _1193;
    wire [191:0] _1202;
    wire [63:0] _1205;
    wire [63:0] data_67;
    wire [63:0] data_68;
    wire [63:0] data_69;
    wire [63:0] data_70;
    wire [5:0] address_70;
    wire _1269;
    wire _1268;
    wire read_enable_58;
    wire _1262 = 1'b0;
    wire _1261 = 1'b0;
    wire _1259 = 1'b0;
    wire _1258 = 1'b0;
    wire _1256 = 1'b0;
    wire _1255 = 1'b0;
    wire _1253 = 1'b0;
    wire _1252 = 1'b0;
    wire _1250 = 1'b0;
    wire _1249 = 1'b0;
    wire _1247 = 1'b0;
    wire _1246 = 1'b0;
    wire _1244 = 1'b0;
    wire _1243 = 1'b0;
    wire _1241 = 1'b0;
    wire _1240 = 1'b0;
    wire _1238 = 1'b0;
    wire _1237 = 1'b0;
    reg _1239;
    reg _1242;
    reg _1245;
    reg _1248;
    reg _1251;
    reg _1254;
    reg _1257;
    reg _1260;
    reg _1263;
    wire _1264;
    wire _1235 = 1'b0;
    wire _1234 = 1'b0;
    wire _1232 = 1'b0;
    wire _1231 = 1'b0;
    wire _1229 = 1'b0;
    wire _1228 = 1'b0;
    wire _1226 = 1'b0;
    wire _1225 = 1'b0;
    wire _1223 = 1'b0;
    wire _1222 = 1'b0;
    wire _1220 = 1'b0;
    wire _1219 = 1'b0;
    wire _1217 = 1'b0;
    wire _1216 = 1'b0;
    wire _1214 = 1'b0;
    wire _1213 = 1'b0;
    wire _1211 = 1'b0;
    wire _1210 = 1'b0;
    reg _1212;
    reg _1215;
    reg _1218;
    reg _1221;
    reg _1224;
    reg _1227;
    reg _1230;
    reg _1233;
    reg _1236;
    wire _1265;
    wire _1266;
    wire write_enable_70;
    wire _1271;
    wire [131:0] _1278;
    wire [63:0] _1279;
    wire _1207 = 1'b0;
    wire _1206 = 1'b0;
    wire _1209;
    wire _47;
    reg PHASE_16;
    wire [63:0] _1291;
    wire [5:0] address_71;
    wire write_enable_71;
    wire [5:0] address_72;
    wire _1466;
    wire read_enable_59;
    wire _1464;
    wire write_enable_72;
    wire _1468;
    wire [131:0] _1473;
    wire [63:0] _1474;
    wire [5:0] _1459 = 6'b000000;
    wire [5:0] address_73;
    wire _1457;
    wire write_enable_73;
    wire [63:0] _1382;
    wire [63:0] _1381;
    wire [63:0] _1383;
    wire [63:0] _1379;
    wire [63:0] _1378;
    wire [63:0] q1_5;
    wire [63:0] _1384;
    wire [5:0] address_74;
    wire write_enable_74 = 1'b0;
    wire _1369;
    wire read_enable_60;
    wire [5:0] address_75;
    wire _1365;
    wire read_enable_61;
    wire _1363;
    wire write_enable_75;
    wire _1367;
    wire [131:0] _1374;
    wire [63:0] _1375;
    wire [63:0] data_71 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_72;
    wire [5:0] _1357 = 6'b000000;
    wire _1355;
    wire _1354;
    wire _1353;
    wire _1352;
    wire _1351;
    wire _1350;
    wire [5:0] _1356;
    wire [5:0] address_76;
    wire write_enable_76 = 1'b0;
    wire _1347;
    wire read_enable_62;
    wire [63:0] data_73;
    wire [63:0] data_74;
    wire _1344;
    wire _1343;
    wire _1342;
    wire _1341;
    wire _1340;
    wire _1339;
    wire [5:0] _1345;
    wire [5:0] address_77;
    wire _1336;
    wire read_enable_63;
    wire _1334;
    wire write_enable_77;
    wire _1338;
    wire [131:0] _1361;
    wire [63:0] _1362;
    wire _1293 = 1'b0;
    wire _1292 = 1'b0;
    wire _1295;
    wire _51;
    reg PHASE_17;
    wire [63:0] _1376;
    wire [5:0] address_78;
    wire _1326;
    wire read_enable_64;
    wire write_enable_78;
    wire _1328;
    wire [5:0] address_79;
    wire _1321;
    wire read_enable_65;
    wire _1319;
    wire write_enable_79;
    wire _1323;
    wire [131:0] _1331;
    wire [63:0] _1332;
    wire [63:0] _1387;
    wire [63:0] data_75;
    wire [63:0] data_76;
    wire [63:0] data_77;
    wire [63:0] data_78;
    wire [5:0] address_80;
    wire _1312;
    wire read_enable_66;
    wire _1309;
    wire _1310;
    wire write_enable_80;
    wire _1314;
    wire [5:0] address_81;
    wire _1305;
    wire read_enable_67;
    wire _1302;
    wire _1303;
    wire write_enable_81;
    wire _1307;
    wire [131:0] _1317;
    wire [63:0] _1318;
    wire _1300 = 1'b0;
    wire _1299 = 1'b0;
    wire _1388;
    wire _53;
    reg PHASE_18;
    wire [63:0] q0_5;
    wire _1297 = 1'b0;
    wire _1296 = 1'b0;
    reg _1298;
    wire [63:0] _1377;
    wire [191:0] _1386;
    wire [63:0] _1389;
    wire [63:0] data_79;
    wire [63:0] data_80;
    wire [63:0] data_81;
    wire [63:0] data_82;
    wire [5:0] address_82;
    wire _1453;
    wire _1452;
    wire read_enable_68;
    wire _1446 = 1'b0;
    wire _1445 = 1'b0;
    wire _1443 = 1'b0;
    wire _1442 = 1'b0;
    wire _1440 = 1'b0;
    wire _1439 = 1'b0;
    wire _1437 = 1'b0;
    wire _1436 = 1'b0;
    wire _1434 = 1'b0;
    wire _1433 = 1'b0;
    wire _1431 = 1'b0;
    wire _1430 = 1'b0;
    wire _1428 = 1'b0;
    wire _1427 = 1'b0;
    wire _1425 = 1'b0;
    wire _1424 = 1'b0;
    wire _1422 = 1'b0;
    wire _1421 = 1'b0;
    reg _1423;
    reg _1426;
    reg _1429;
    reg _1432;
    reg _1435;
    reg _1438;
    reg _1441;
    reg _1444;
    reg _1447;
    wire _1448;
    wire _1419 = 1'b0;
    wire _1418 = 1'b0;
    wire _1416 = 1'b0;
    wire _1415 = 1'b0;
    wire _1413 = 1'b0;
    wire _1412 = 1'b0;
    wire _1410 = 1'b0;
    wire _1409 = 1'b0;
    wire _1407 = 1'b0;
    wire _1406 = 1'b0;
    wire _1404 = 1'b0;
    wire _1403 = 1'b0;
    wire _1401 = 1'b0;
    wire _1400 = 1'b0;
    wire _1398 = 1'b0;
    wire _1397 = 1'b0;
    wire _1395 = 1'b0;
    wire _1394 = 1'b0;
    reg _1396;
    reg _1399;
    reg _1402;
    reg _1405;
    reg _1408;
    reg _1411;
    reg _1414;
    reg _1417;
    reg _1420;
    wire _1449;
    wire _1450;
    wire write_enable_82;
    wire _1455;
    wire [131:0] _1462;
    wire [63:0] _1463;
    wire _1391 = 1'b0;
    wire _1390 = 1'b0;
    wire _1393;
    wire _55;
    reg PHASE_19;
    wire [63:0] _1475;
    wire [5:0] address_83;
    wire write_enable_83;
    wire [5:0] address_84;
    wire _1650;
    wire read_enable_69;
    wire _1648;
    wire write_enable_84;
    wire _1652;
    wire [131:0] _1657;
    wire [63:0] _1658;
    wire [5:0] _1643 = 6'b000000;
    wire [5:0] address_85;
    wire _1641;
    wire write_enable_85;
    wire [3:0] _280;
    wire _279;
    wire _277;
    wire [63:0] _276;
    wire [63:0] _275;
    wire [63:0] _274;
    wire [63:0] _273;
    wire [63:0] _272;
    wire [63:0] _271;
    wire [63:0] _270;
    wire [63:0] _1566;
    wire [63:0] _1565;
    wire [63:0] _1567;
    wire [63:0] _1563;
    wire [63:0] _1562;
    wire [63:0] q1_6;
    wire [63:0] _1568;
    wire [5:0] address_86;
    wire write_enable_86 = 1'b0;
    wire _1553;
    wire read_enable_70;
    wire [5:0] address_87;
    wire _1549;
    wire read_enable_71;
    wire _1547;
    wire write_enable_87;
    wire _1551;
    wire [131:0] _1558;
    wire [63:0] _1559;
    wire [63:0] data_83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_84;
    wire [5:0] _1541 = 6'b000000;
    wire _1539;
    wire _1538;
    wire _1537;
    wire _1536;
    wire _1535;
    wire _1534;
    wire [5:0] _1540;
    wire [5:0] address_88;
    wire write_enable_88 = 1'b0;
    wire _1531;
    wire read_enable_72;
    wire [63:0] data_85;
    wire [63:0] data_86;
    wire [5:0] _60;
    wire _1528;
    wire _1527;
    wire _1526;
    wire _1525;
    wire _1524;
    wire _1523;
    wire [5:0] _1529;
    wire [5:0] address_89;
    wire _1520;
    wire read_enable_73;
    wire [7:0] _62;
    wire _1518;
    wire write_enable_89;
    wire _1522;
    wire [131:0] _1545;
    wire [63:0] _1546;
    wire _1477 = 1'b0;
    wire _1476 = 1'b0;
    wire _1479;
    wire _63;
    reg PHASE_20;
    wire [63:0] _1560;
    wire [5:0] address_90;
    wire _1510;
    wire read_enable_74;
    wire write_enable_90;
    wire _1512;
    wire [5:0] address_91;
    wire _1505;
    wire read_enable_75;
    wire _1503;
    wire write_enable_91;
    wire _1507;
    wire [131:0] _1515;
    wire [63:0] _1516;
    wire [63:0] _1571;
    wire [63:0] data_87;
    wire [63:0] data_88;
    wire [63:0] data_89;
    wire [63:0] data_90;
    wire [5:0] _198 = 6'b000000;
    wire [5:0] _197 = 6'b000000;
    wire [5:0] _195 = 6'b000000;
    wire [5:0] _194 = 6'b000000;
    wire [5:0] _192 = 6'b000000;
    wire [5:0] _191 = 6'b000000;
    wire [5:0] _189 = 6'b000000;
    wire [5:0] _188 = 6'b000000;
    wire [5:0] _186 = 6'b000000;
    wire [5:0] _185 = 6'b000000;
    wire [5:0] _183 = 6'b000000;
    wire [5:0] _182 = 6'b000000;
    wire [5:0] _180 = 6'b000000;
    wire [5:0] _179 = 6'b000000;
    wire [5:0] _177 = 6'b000000;
    wire [5:0] _176 = 6'b000000;
    wire [5:0] _174 = 6'b000000;
    wire [5:0] _173 = 6'b000000;
    reg [5:0] _175;
    reg [5:0] _178;
    reg [5:0] _181;
    reg [5:0] _184;
    reg [5:0] _187;
    reg [5:0] _190;
    reg [5:0] _193;
    reg [5:0] _196;
    reg [5:0] _199;
    wire [5:0] _172;
    wire [5:0] address_92;
    wire _1496;
    wire read_enable_76;
    wire _1493;
    wire _1494;
    wire write_enable_92;
    wire _1498;
    wire [5:0] address_93;
    wire _1489;
    wire read_enable_77;
    wire _1486;
    wire _1487;
    wire write_enable_93;
    wire _1491;
    wire [131:0] _1501;
    wire [63:0] _1502;
    wire _99;
    wire _1484 = 1'b0;
    wire _1483 = 1'b0;
    wire _1572;
    wire _65;
    reg PHASE_21;
    wire [63:0] q0_6;
    wire _1481 = 1'b0;
    wire _1480 = 1'b0;
    wire _92;
    reg _1482;
    wire [63:0] _1561;
    wire [191:0] _1570;
    wire [63:0] _1573;
    wire [63:0] data_91;
    wire [63:0] data_92;
    wire [63:0] data_93;
    wire [63:0] data_94;
    wire [5:0] _163 = 6'b000000;
    wire [5:0] _162 = 6'b000000;
    wire [5:0] _160 = 6'b000000;
    wire [5:0] _159 = 6'b000000;
    wire [5:0] _157 = 6'b000000;
    wire [5:0] _156 = 6'b000000;
    wire [5:0] _154 = 6'b000000;
    wire [5:0] _153 = 6'b000000;
    wire [5:0] _151 = 6'b000000;
    wire [5:0] _150 = 6'b000000;
    wire [5:0] _148 = 6'b000000;
    wire [5:0] _147 = 6'b000000;
    wire [5:0] _145 = 6'b000000;
    wire [5:0] _144 = 6'b000000;
    wire [5:0] _142 = 6'b000000;
    wire [5:0] _141 = 6'b000000;
    wire [5:0] _139 = 6'b000000;
    wire [5:0] _138 = 6'b000000;
    wire [5:0] _137;
    reg [5:0] _140;
    reg [5:0] _143;
    reg [5:0] _146;
    reg [5:0] _149;
    reg [5:0] _152;
    reg [5:0] _155;
    reg [5:0] _158;
    reg [5:0] _161;
    reg [5:0] _164;
    wire [5:0] _68;
    wire [5:0] address_94;
    wire _1637;
    wire [7:0] _70;
    wire _1636;
    wire read_enable_78;
    wire _1630 = 1'b0;
    wire _1629 = 1'b0;
    wire _1627 = 1'b0;
    wire _1626 = 1'b0;
    wire _1624 = 1'b0;
    wire _1623 = 1'b0;
    wire _1621 = 1'b0;
    wire _1620 = 1'b0;
    wire _1618 = 1'b0;
    wire _1617 = 1'b0;
    wire _1615 = 1'b0;
    wire _1614 = 1'b0;
    wire _1612 = 1'b0;
    wire _1611 = 1'b0;
    wire _1609 = 1'b0;
    wire _1608 = 1'b0;
    wire _1606 = 1'b0;
    wire _1605 = 1'b0;
    wire _278;
    reg _1607;
    reg _1610;
    reg _1613;
    reg _1616;
    reg _1619;
    reg _1622;
    reg _1625;
    reg _1628;
    reg _1631;
    wire _1632;
    wire _1603 = 1'b0;
    wire _1602 = 1'b0;
    wire _1600 = 1'b0;
    wire _1599 = 1'b0;
    wire _1597 = 1'b0;
    wire _1596 = 1'b0;
    wire _1594 = 1'b0;
    wire _1593 = 1'b0;
    wire _1591 = 1'b0;
    wire _1590 = 1'b0;
    wire _1588 = 1'b0;
    wire _1587 = 1'b0;
    wire _1585 = 1'b0;
    wire _1584 = 1'b0;
    wire _1582 = 1'b0;
    wire _1581 = 1'b0;
    wire _1579 = 1'b0;
    wire _1578 = 1'b0;
    wire _130;
    reg _1580;
    reg _1583;
    reg _1586;
    reg _1589;
    reg _1592;
    reg _1595;
    reg _1598;
    reg _1601;
    reg _1604;
    wire _1633;
    wire _128 = 1'b0;
    wire _127 = 1'b0;
    wire _125 = 1'b0;
    wire _124 = 1'b0;
    wire _122 = 1'b0;
    wire _121 = 1'b0;
    wire _119 = 1'b0;
    wire _118 = 1'b0;
    wire _116 = 1'b0;
    wire _115 = 1'b0;
    wire _113 = 1'b0;
    wire _112 = 1'b0;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire vdd = 1'b1;
    wire _104 = 1'b0;
    wire _103 = 1'b0;
    wire _102;
    reg _105;
    reg _108;
    reg _111;
    reg _114;
    reg _117;
    reg _120;
    reg _123;
    reg _126;
    reg _129;
    wire _1634;
    wire write_enable_94;
    wire _1639;
    wire gnd = 1'b0;
    wire [131:0] _1646;
    wire [63:0] _1647;
    wire _72;
    wire _1575 = 1'b0;
    wire _1574 = 1'b0;
    wire _1577;
    wire _73;
    reg PHASE_22;
    wire [63:0] _1659;
    wire _76;
    wire _78;
    wire _80;
    wire _82;
    wire _84;
    wire [492:0] _91;
    wire _1660;

    /* logic */
    assign address = _360 ? _199 : _355;
    assign write_enable = _353 & _360;
    assign address_0 = _360 ? _164 : _68;
    assign _362 = ~ _360;
    assign read_enable = _348 & _362;
    assign _360 = ~ PHASE_1;
    assign write_enable_0 = _346 & _360;
    assign _364 = write_enable_0 | read_enable;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_364), .regcea(vdd), .wea(write_enable_0), .addra(address_0), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable), .regceb(vdd), .web(write_enable), .addrb(address), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_369[131:131]), .sbiterrb(_369[130:130]), .doutb(_369[129:66]), .dbiterra(_369[65:65]), .sbiterra(_369[64:64]), .douta(_369[63:0]) );
    assign _370 = _369[63:0];
    assign address_1 = PHASE_1 ? _199 : _355;
    assign _353 = _129 & _316;
    assign write_enable_1 = _353 & PHASE_1;
    assign _267 = _259[129:66];
    assign _266 = _246[129:66];
    assign _268 = PHASE ? _267 : _266;
    assign _264 = _216[129:66];
    assign _263 = _202[129:66];
    assign q1 = PHASE_0 ? _264 : _263;
    assign _269 = _96 ? _268 : q1;
    assign address_2 = _248 ? _242 : _241;
    assign _254 = ~ _248;
    assign read_enable_0 = _102 & _254;
    assign address_3 = _248 ? _60 : _230;
    assign _250 = ~ _248;
    assign read_enable_1 = _102 & _250;
    assign _248 = ~ PHASE;
    assign write_enable_3 = _219 & _248;
    assign _252 = write_enable_3 | read_enable_1;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_0
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_252), .regcea(vdd), .wea(write_enable_3), .addra(address_3), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_0), .regceb(vdd), .web(write_enable_2), .addrb(address_2), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_259[131:131]), .sbiterrb(_259[130:130]), .doutb(_259[129:66]), .dbiterra(_259[65:65]), .sbiterra(_259[64:64]), .douta(_259[63:0]) );
    assign _260 = _259[63:0];
    assign _240 = _172[5:5];
    assign _239 = _172[4:4];
    assign _238 = _172[3:3];
    assign _237 = _172[2:2];
    assign _236 = _172[1:1];
    assign _235 = _172[0:0];
    assign _241 = { _235, _236, _237, _238, _239, _240 };
    assign address_4 = PHASE ? _242 : _241;
    assign _232 = ~ PHASE;
    assign read_enable_2 = _102 & _232;
    assign data_1 = wr_d7;
    assign _229 = _137[5:5];
    assign _228 = _137[4:4];
    assign _227 = _137[3:3];
    assign _226 = _137[2:2];
    assign _225 = _137[1:1];
    assign _224 = _137[0:0];
    assign _230 = { _224, _225, _226, _227, _228, _229 };
    assign address_5 = PHASE ? _60 : _230;
    assign _221 = ~ PHASE;
    assign read_enable_3 = _102 & _221;
    assign _219 = _62[7:7];
    assign write_enable_5 = _219 & PHASE;
    assign _223 = write_enable_5 | read_enable_3;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_1
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_223), .regcea(vdd), .wea(write_enable_5), .addra(address_5), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_2), .regceb(vdd), .web(write_enable_4), .addrb(address_4), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_246[131:131]), .sbiterrb(_246[130:130]), .doutb(_246[129:66]), .dbiterra(_246[65:65]), .sbiterra(_246[64:64]), .douta(_246[63:0]) );
    assign _247 = _246[63:0];
    assign _89 = ~ PHASE;
    assign _3 = _89;
    always @(posedge _84) begin
        if (_82)
            PHASE <= _87;
        else
            if (_72)
                PHASE <= _3;
    end
    assign _261 = PHASE ? _260 : _247;
    assign address_6 = _204 ? _199 : _172;
    assign _211 = ~ _204;
    assign read_enable_4 = _102 & _211;
    assign write_enable_6 = _167 & _204;
    assign _213 = write_enable_6 | read_enable_4;
    assign address_7 = _204 ? _164 : _137;
    assign _206 = ~ _204;
    assign read_enable_5 = _102 & _206;
    assign _204 = ~ PHASE_0;
    assign write_enable_7 = _132 & _204;
    assign _208 = write_enable_7 | read_enable_5;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_2
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_208), .regcea(vdd), .wea(write_enable_7), .addra(address_7), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_213), .regceb(vdd), .web(write_enable_6), .addrb(address_6), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_216[131:131]), .sbiterrb(_216[130:130]), .doutb(_216[129:66]), .dbiterra(_216[65:65]), .sbiterra(_216[64:64]), .douta(_216[63:0]) );
    assign _217 = _216[63:0];
    assign _283 = _282[127:64];
    assign data_3 = _283;
    assign address_8 = PHASE_0 ? _199 : _172;
    assign _169 = ~ PHASE_0;
    assign read_enable_6 = _102 & _169;
    assign _166 = ~ _130;
    assign _167 = _129 & _166;
    assign write_enable_8 = _167 & PHASE_0;
    assign _171 = write_enable_8 | read_enable_6;
    assign address_9 = PHASE_0 ? _164 : _137;
    assign _134 = ~ PHASE_0;
    assign read_enable_7 = _102 & _134;
    assign _131 = ~ _130;
    assign _132 = _129 & _131;
    assign write_enable_9 = _132 & PHASE_0;
    assign _136 = write_enable_9 | read_enable_7;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_3
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_136), .regcea(vdd), .wea(write_enable_9), .addra(address_9), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_171), .regceb(vdd), .web(write_enable_8), .addrb(address_8), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_202[131:131]), .sbiterrb(_202[130:130]), .doutb(_202[129:66]), .dbiterra(_202[65:65]), .sbiterra(_202[64:64]), .douta(_202[63:0]) );
    assign _203 = _202[63:0];
    assign _284 = ~ PHASE_0;
    assign _5 = _284;
    always @(posedge _84) begin
        if (_82)
            PHASE_0 <= _98;
        else
            if (_99)
                PHASE_0 <= _5;
    end
    assign q0 = PHASE_0 ? _217 : _203;
    always @(posedge _84) begin
        if (_82)
            _96 <= _94;
        else
            _96 <= _92;
    end
    assign _262 = _96 ? _261 : q0;
    dp_22
        dp_6
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_262), .d2(_269), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_282[191:128]), .q2(_282[127:64]), .q1(_282[63:0]) );
    assign _285 = _282[63:0];
    assign data_7 = _285;
    assign address_10 = PHASE_1 ? _164 : _68;
    assign _349 = ~ PHASE_1;
    assign _348 = _70[7:7];
    assign read_enable_8 = _348 & _349;
    always @(posedge _84) begin
        if (_82)
            _319 <= _318;
        else
            _319 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _322 <= _321;
        else
            _322 <= _319;
    end
    always @(posedge _84) begin
        if (_82)
            _325 <= _324;
        else
            _325 <= _322;
    end
    always @(posedge _84) begin
        if (_82)
            _328 <= _327;
        else
            _328 <= _325;
    end
    always @(posedge _84) begin
        if (_82)
            _331 <= _330;
        else
            _331 <= _328;
    end
    always @(posedge _84) begin
        if (_82)
            _334 <= _333;
        else
            _334 <= _331;
    end
    always @(posedge _84) begin
        if (_82)
            _337 <= _336;
        else
            _337 <= _334;
    end
    always @(posedge _84) begin
        if (_82)
            _340 <= _339;
        else
            _340 <= _337;
    end
    always @(posedge _84) begin
        if (_82)
            _343 <= _342;
        else
            _343 <= _340;
    end
    assign _344 = ~ _343;
    always @(posedge _84) begin
        if (_82)
            _292 <= _291;
        else
            _292 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _295 <= _294;
        else
            _295 <= _292;
    end
    always @(posedge _84) begin
        if (_82)
            _298 <= _297;
        else
            _298 <= _295;
    end
    always @(posedge _84) begin
        if (_82)
            _301 <= _300;
        else
            _301 <= _298;
    end
    always @(posedge _84) begin
        if (_82)
            _304 <= _303;
        else
            _304 <= _301;
    end
    always @(posedge _84) begin
        if (_82)
            _307 <= _306;
        else
            _307 <= _304;
    end
    always @(posedge _84) begin
        if (_82)
            _310 <= _309;
        else
            _310 <= _307;
    end
    always @(posedge _84) begin
        if (_82)
            _313 <= _312;
        else
            _313 <= _310;
    end
    always @(posedge _84) begin
        if (_82)
            _316 <= _315;
        else
            _316 <= _313;
    end
    assign _345 = _316 & _344;
    assign _346 = _129 & _345;
    assign write_enable_10 = _346 & PHASE_1;
    assign _351 = write_enable_10 | read_enable_8;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_4
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_351), .regcea(vdd), .wea(write_enable_10), .addra(address_10), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_1), .regceb(vdd), .web(write_enable_1), .addrb(address_1), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_358[131:131]), .sbiterrb(_358[130:130]), .doutb(_358[129:66]), .dbiterra(_358[65:65]), .sbiterra(_358[64:64]), .douta(_358[63:0]) );
    assign _359 = _358[63:0];
    assign _289 = ~ PHASE_1;
    assign _7 = _289;
    always @(posedge _84) begin
        if (_82)
            PHASE_1 <= _287;
        else
            if (_72)
                PHASE_1 <= _7;
    end
    assign _371 = PHASE_1 ? _370 : _359;
    assign address_11 = _544 ? _199 : _539;
    assign write_enable_11 = _537 & _544;
    assign address_12 = _544 ? _164 : _68;
    assign _546 = ~ _544;
    assign read_enable_9 = _532 & _546;
    assign _544 = ~ PHASE_4;
    assign write_enable_12 = _530 & _544;
    assign _548 = write_enable_12 | read_enable_9;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_5
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_548), .regcea(vdd), .wea(write_enable_12), .addra(address_12), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_11), .regceb(vdd), .web(write_enable_11), .addrb(address_11), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_553[131:131]), .sbiterrb(_553[130:130]), .doutb(_553[129:66]), .dbiterra(_553[65:65]), .sbiterra(_553[64:64]), .douta(_553[63:0]) );
    assign _554 = _553[63:0];
    assign address_13 = PHASE_4 ? _199 : _539;
    assign _537 = _129 & _500;
    assign write_enable_13 = _537 & PHASE_4;
    assign _462 = _454[129:66];
    assign _461 = _441[129:66];
    assign _463 = PHASE_2 ? _462 : _461;
    assign _459 = _411[129:66];
    assign _458 = _397[129:66];
    assign q1_0 = PHASE_3 ? _459 : _458;
    assign _464 = _378 ? _463 : q1_0;
    assign address_14 = _443 ? _437 : _436;
    assign _449 = ~ _443;
    assign read_enable_10 = _102 & _449;
    assign address_15 = _443 ? _60 : _425;
    assign _445 = ~ _443;
    assign read_enable_11 = _102 & _445;
    assign _443 = ~ PHASE_2;
    assign write_enable_15 = _414 & _443;
    assign _447 = write_enable_15 | read_enable_11;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_6
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_447), .regcea(vdd), .wea(write_enable_15), .addra(address_15), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_10), .regceb(vdd), .web(write_enable_14), .addrb(address_14), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_454[131:131]), .sbiterrb(_454[130:130]), .doutb(_454[129:66]), .dbiterra(_454[65:65]), .sbiterra(_454[64:64]), .douta(_454[63:0]) );
    assign _455 = _454[63:0];
    assign _435 = _172[5:5];
    assign _434 = _172[4:4];
    assign _433 = _172[3:3];
    assign _432 = _172[2:2];
    assign _431 = _172[1:1];
    assign _430 = _172[0:0];
    assign _436 = { _430, _431, _432, _433, _434, _435 };
    assign address_16 = PHASE_2 ? _437 : _436;
    assign _427 = ~ PHASE_2;
    assign read_enable_12 = _102 & _427;
    assign data_13 = wr_d6;
    assign _424 = _137[5:5];
    assign _423 = _137[4:4];
    assign _422 = _137[3:3];
    assign _421 = _137[2:2];
    assign _420 = _137[1:1];
    assign _419 = _137[0:0];
    assign _425 = { _419, _420, _421, _422, _423, _424 };
    assign address_17 = PHASE_2 ? _60 : _425;
    assign _416 = ~ PHASE_2;
    assign read_enable_13 = _102 & _416;
    assign _414 = _62[6:6];
    assign write_enable_17 = _414 & PHASE_2;
    assign _418 = write_enable_17 | read_enable_13;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_7
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_418), .regcea(vdd), .wea(write_enable_17), .addra(address_17), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_12), .regceb(vdd), .web(write_enable_16), .addrb(address_16), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_441[131:131]), .sbiterrb(_441[130:130]), .doutb(_441[129:66]), .dbiterra(_441[65:65]), .sbiterra(_441[64:64]), .douta(_441[63:0]) );
    assign _442 = _441[63:0];
    assign _375 = ~ PHASE_2;
    assign _11 = _375;
    always @(posedge _84) begin
        if (_82)
            PHASE_2 <= _373;
        else
            if (_72)
                PHASE_2 <= _11;
    end
    assign _456 = PHASE_2 ? _455 : _442;
    assign address_18 = _399 ? _199 : _172;
    assign _406 = ~ _399;
    assign read_enable_14 = _102 & _406;
    assign write_enable_18 = _390 & _399;
    assign _408 = write_enable_18 | read_enable_14;
    assign address_19 = _399 ? _164 : _137;
    assign _401 = ~ _399;
    assign read_enable_15 = _102 & _401;
    assign _399 = ~ PHASE_3;
    assign write_enable_19 = _383 & _399;
    assign _403 = write_enable_19 | read_enable_15;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_8
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_403), .regcea(vdd), .wea(write_enable_19), .addra(address_19), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_408), .regceb(vdd), .web(write_enable_18), .addrb(address_18), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_411[131:131]), .sbiterrb(_411[130:130]), .doutb(_411[129:66]), .dbiterra(_411[65:65]), .sbiterra(_411[64:64]), .douta(_411[63:0]) );
    assign _412 = _411[63:0];
    assign _467 = _466[127:64];
    assign data_15 = _467;
    assign address_20 = PHASE_3 ? _199 : _172;
    assign _392 = ~ PHASE_3;
    assign read_enable_16 = _102 & _392;
    assign _389 = ~ _130;
    assign _390 = _129 & _389;
    assign write_enable_20 = _390 & PHASE_3;
    assign _394 = write_enable_20 | read_enable_16;
    assign address_21 = PHASE_3 ? _164 : _137;
    assign _385 = ~ PHASE_3;
    assign read_enable_17 = _102 & _385;
    assign _382 = ~ _130;
    assign _383 = _129 & _382;
    assign write_enable_21 = _383 & PHASE_3;
    assign _387 = write_enable_21 | read_enable_17;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_9
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_387), .regcea(vdd), .wea(write_enable_21), .addra(address_21), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_394), .regceb(vdd), .web(write_enable_20), .addrb(address_20), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_397[131:131]), .sbiterrb(_397[130:130]), .doutb(_397[129:66]), .dbiterra(_397[65:65]), .sbiterra(_397[64:64]), .douta(_397[63:0]) );
    assign _398 = _397[63:0];
    assign _468 = ~ PHASE_3;
    assign _13 = _468;
    always @(posedge _84) begin
        if (_82)
            PHASE_3 <= _380;
        else
            if (_99)
                PHASE_3 <= _13;
    end
    assign q0_0 = PHASE_3 ? _412 : _398;
    always @(posedge _84) begin
        if (_82)
            _378 <= _377;
        else
            _378 <= _92;
    end
    assign _457 = _378 ? _456 : q0_0;
    dp_21
        dp_5
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_457), .d2(_464), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_466[191:128]), .q2(_466[127:64]), .q1(_466[63:0]) );
    assign _469 = _466[63:0];
    assign data_19 = _469;
    assign address_22 = PHASE_4 ? _164 : _68;
    assign _533 = ~ PHASE_4;
    assign _532 = _70[6:6];
    assign read_enable_18 = _532 & _533;
    always @(posedge _84) begin
        if (_82)
            _503 <= _502;
        else
            _503 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _506 <= _505;
        else
            _506 <= _503;
    end
    always @(posedge _84) begin
        if (_82)
            _509 <= _508;
        else
            _509 <= _506;
    end
    always @(posedge _84) begin
        if (_82)
            _512 <= _511;
        else
            _512 <= _509;
    end
    always @(posedge _84) begin
        if (_82)
            _515 <= _514;
        else
            _515 <= _512;
    end
    always @(posedge _84) begin
        if (_82)
            _518 <= _517;
        else
            _518 <= _515;
    end
    always @(posedge _84) begin
        if (_82)
            _521 <= _520;
        else
            _521 <= _518;
    end
    always @(posedge _84) begin
        if (_82)
            _524 <= _523;
        else
            _524 <= _521;
    end
    always @(posedge _84) begin
        if (_82)
            _527 <= _526;
        else
            _527 <= _524;
    end
    assign _528 = ~ _527;
    always @(posedge _84) begin
        if (_82)
            _476 <= _475;
        else
            _476 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _479 <= _478;
        else
            _479 <= _476;
    end
    always @(posedge _84) begin
        if (_82)
            _482 <= _481;
        else
            _482 <= _479;
    end
    always @(posedge _84) begin
        if (_82)
            _485 <= _484;
        else
            _485 <= _482;
    end
    always @(posedge _84) begin
        if (_82)
            _488 <= _487;
        else
            _488 <= _485;
    end
    always @(posedge _84) begin
        if (_82)
            _491 <= _490;
        else
            _491 <= _488;
    end
    always @(posedge _84) begin
        if (_82)
            _494 <= _493;
        else
            _494 <= _491;
    end
    always @(posedge _84) begin
        if (_82)
            _497 <= _496;
        else
            _497 <= _494;
    end
    always @(posedge _84) begin
        if (_82)
            _500 <= _499;
        else
            _500 <= _497;
    end
    assign _529 = _500 & _528;
    assign _530 = _129 & _529;
    assign write_enable_22 = _530 & PHASE_4;
    assign _535 = write_enable_22 | read_enable_18;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_10
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_535), .regcea(vdd), .wea(write_enable_22), .addra(address_22), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_13), .regceb(vdd), .web(write_enable_13), .addrb(address_13), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_542[131:131]), .sbiterrb(_542[130:130]), .doutb(_542[129:66]), .dbiterra(_542[65:65]), .sbiterra(_542[64:64]), .douta(_542[63:0]) );
    assign _543 = _542[63:0];
    assign _473 = ~ PHASE_4;
    assign _15 = _473;
    always @(posedge _84) begin
        if (_82)
            PHASE_4 <= _471;
        else
            if (_72)
                PHASE_4 <= _15;
    end
    assign _555 = PHASE_4 ? _554 : _543;
    assign address_23 = _728 ? _199 : _723;
    assign write_enable_23 = _721 & _728;
    assign address_24 = _728 ? _164 : _68;
    assign _730 = ~ _728;
    assign read_enable_19 = _716 & _730;
    assign _728 = ~ PHASE_7;
    assign write_enable_24 = _714 & _728;
    assign _732 = write_enable_24 | read_enable_19;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_11
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_732), .regcea(vdd), .wea(write_enable_24), .addra(address_24), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_23), .regceb(vdd), .web(write_enable_23), .addrb(address_23), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_737[131:131]), .sbiterrb(_737[130:130]), .doutb(_737[129:66]), .dbiterra(_737[65:65]), .sbiterra(_737[64:64]), .douta(_737[63:0]) );
    assign _738 = _737[63:0];
    assign address_25 = PHASE_7 ? _199 : _723;
    assign _721 = _129 & _684;
    assign write_enable_25 = _721 & PHASE_7;
    assign _646 = _638[129:66];
    assign _645 = _625[129:66];
    assign _647 = PHASE_5 ? _646 : _645;
    assign _643 = _595[129:66];
    assign _642 = _581[129:66];
    assign q1_1 = PHASE_6 ? _643 : _642;
    assign _648 = _562 ? _647 : q1_1;
    assign address_26 = _627 ? _621 : _620;
    assign _633 = ~ _627;
    assign read_enable_20 = _102 & _633;
    assign address_27 = _627 ? _60 : _609;
    assign _629 = ~ _627;
    assign read_enable_21 = _102 & _629;
    assign _627 = ~ PHASE_5;
    assign write_enable_27 = _598 & _627;
    assign _631 = write_enable_27 | read_enable_21;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_12
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_631), .regcea(vdd), .wea(write_enable_27), .addra(address_27), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_20), .regceb(vdd), .web(write_enable_26), .addrb(address_26), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_638[131:131]), .sbiterrb(_638[130:130]), .doutb(_638[129:66]), .dbiterra(_638[65:65]), .sbiterra(_638[64:64]), .douta(_638[63:0]) );
    assign _639 = _638[63:0];
    assign _619 = _172[5:5];
    assign _618 = _172[4:4];
    assign _617 = _172[3:3];
    assign _616 = _172[2:2];
    assign _615 = _172[1:1];
    assign _614 = _172[0:0];
    assign _620 = { _614, _615, _616, _617, _618, _619 };
    assign address_28 = PHASE_5 ? _621 : _620;
    assign _611 = ~ PHASE_5;
    assign read_enable_22 = _102 & _611;
    assign data_25 = wr_d5;
    assign _608 = _137[5:5];
    assign _607 = _137[4:4];
    assign _606 = _137[3:3];
    assign _605 = _137[2:2];
    assign _604 = _137[1:1];
    assign _603 = _137[0:0];
    assign _609 = { _603, _604, _605, _606, _607, _608 };
    assign address_29 = PHASE_5 ? _60 : _609;
    assign _600 = ~ PHASE_5;
    assign read_enable_23 = _102 & _600;
    assign _598 = _62[5:5];
    assign write_enable_29 = _598 & PHASE_5;
    assign _602 = write_enable_29 | read_enable_23;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_13
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_602), .regcea(vdd), .wea(write_enable_29), .addra(address_29), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_22), .regceb(vdd), .web(write_enable_28), .addrb(address_28), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_625[131:131]), .sbiterrb(_625[130:130]), .doutb(_625[129:66]), .dbiterra(_625[65:65]), .sbiterra(_625[64:64]), .douta(_625[63:0]) );
    assign _626 = _625[63:0];
    assign _559 = ~ PHASE_5;
    assign _19 = _559;
    always @(posedge _84) begin
        if (_82)
            PHASE_5 <= _557;
        else
            if (_72)
                PHASE_5 <= _19;
    end
    assign _640 = PHASE_5 ? _639 : _626;
    assign address_30 = _583 ? _199 : _172;
    assign _590 = ~ _583;
    assign read_enable_24 = _102 & _590;
    assign write_enable_30 = _574 & _583;
    assign _592 = write_enable_30 | read_enable_24;
    assign address_31 = _583 ? _164 : _137;
    assign _585 = ~ _583;
    assign read_enable_25 = _102 & _585;
    assign _583 = ~ PHASE_6;
    assign write_enable_31 = _567 & _583;
    assign _587 = write_enable_31 | read_enable_25;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_14
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_587), .regcea(vdd), .wea(write_enable_31), .addra(address_31), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_592), .regceb(vdd), .web(write_enable_30), .addrb(address_30), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_595[131:131]), .sbiterrb(_595[130:130]), .doutb(_595[129:66]), .dbiterra(_595[65:65]), .sbiterra(_595[64:64]), .douta(_595[63:0]) );
    assign _596 = _595[63:0];
    assign _651 = _650[127:64];
    assign data_27 = _651;
    assign address_32 = PHASE_6 ? _199 : _172;
    assign _576 = ~ PHASE_6;
    assign read_enable_26 = _102 & _576;
    assign _573 = ~ _130;
    assign _574 = _129 & _573;
    assign write_enable_32 = _574 & PHASE_6;
    assign _578 = write_enable_32 | read_enable_26;
    assign address_33 = PHASE_6 ? _164 : _137;
    assign _569 = ~ PHASE_6;
    assign read_enable_27 = _102 & _569;
    assign _566 = ~ _130;
    assign _567 = _129 & _566;
    assign write_enable_33 = _567 & PHASE_6;
    assign _571 = write_enable_33 | read_enable_27;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_15
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_571), .regcea(vdd), .wea(write_enable_33), .addra(address_33), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_578), .regceb(vdd), .web(write_enable_32), .addrb(address_32), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_581[131:131]), .sbiterrb(_581[130:130]), .doutb(_581[129:66]), .dbiterra(_581[65:65]), .sbiterra(_581[64:64]), .douta(_581[63:0]) );
    assign _582 = _581[63:0];
    assign _652 = ~ PHASE_6;
    assign _21 = _652;
    always @(posedge _84) begin
        if (_82)
            PHASE_6 <= _564;
        else
            if (_99)
                PHASE_6 <= _21;
    end
    assign q0_1 = PHASE_6 ? _596 : _582;
    always @(posedge _84) begin
        if (_82)
            _562 <= _561;
        else
            _562 <= _92;
    end
    assign _641 = _562 ? _640 : q0_1;
    dp_20
        dp_4
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_641), .d2(_648), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_650[191:128]), .q2(_650[127:64]), .q1(_650[63:0]) );
    assign _653 = _650[63:0];
    assign data_31 = _653;
    assign address_34 = PHASE_7 ? _164 : _68;
    assign _717 = ~ PHASE_7;
    assign _716 = _70[5:5];
    assign read_enable_28 = _716 & _717;
    always @(posedge _84) begin
        if (_82)
            _687 <= _686;
        else
            _687 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _690 <= _689;
        else
            _690 <= _687;
    end
    always @(posedge _84) begin
        if (_82)
            _693 <= _692;
        else
            _693 <= _690;
    end
    always @(posedge _84) begin
        if (_82)
            _696 <= _695;
        else
            _696 <= _693;
    end
    always @(posedge _84) begin
        if (_82)
            _699 <= _698;
        else
            _699 <= _696;
    end
    always @(posedge _84) begin
        if (_82)
            _702 <= _701;
        else
            _702 <= _699;
    end
    always @(posedge _84) begin
        if (_82)
            _705 <= _704;
        else
            _705 <= _702;
    end
    always @(posedge _84) begin
        if (_82)
            _708 <= _707;
        else
            _708 <= _705;
    end
    always @(posedge _84) begin
        if (_82)
            _711 <= _710;
        else
            _711 <= _708;
    end
    assign _712 = ~ _711;
    always @(posedge _84) begin
        if (_82)
            _660 <= _659;
        else
            _660 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _663 <= _662;
        else
            _663 <= _660;
    end
    always @(posedge _84) begin
        if (_82)
            _666 <= _665;
        else
            _666 <= _663;
    end
    always @(posedge _84) begin
        if (_82)
            _669 <= _668;
        else
            _669 <= _666;
    end
    always @(posedge _84) begin
        if (_82)
            _672 <= _671;
        else
            _672 <= _669;
    end
    always @(posedge _84) begin
        if (_82)
            _675 <= _674;
        else
            _675 <= _672;
    end
    always @(posedge _84) begin
        if (_82)
            _678 <= _677;
        else
            _678 <= _675;
    end
    always @(posedge _84) begin
        if (_82)
            _681 <= _680;
        else
            _681 <= _678;
    end
    always @(posedge _84) begin
        if (_82)
            _684 <= _683;
        else
            _684 <= _681;
    end
    assign _713 = _684 & _712;
    assign _714 = _129 & _713;
    assign write_enable_34 = _714 & PHASE_7;
    assign _719 = write_enable_34 | read_enable_28;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_16
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_719), .regcea(vdd), .wea(write_enable_34), .addra(address_34), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_25), .regceb(vdd), .web(write_enable_25), .addrb(address_25), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_726[131:131]), .sbiterrb(_726[130:130]), .doutb(_726[129:66]), .dbiterra(_726[65:65]), .sbiterra(_726[64:64]), .douta(_726[63:0]) );
    assign _727 = _726[63:0];
    assign _657 = ~ PHASE_7;
    assign _23 = _657;
    always @(posedge _84) begin
        if (_82)
            PHASE_7 <= _655;
        else
            if (_72)
                PHASE_7 <= _23;
    end
    assign _739 = PHASE_7 ? _738 : _727;
    assign address_35 = _912 ? _199 : _907;
    assign write_enable_35 = _905 & _912;
    assign address_36 = _912 ? _164 : _68;
    assign _914 = ~ _912;
    assign read_enable_29 = _900 & _914;
    assign _912 = ~ PHASE_10;
    assign write_enable_36 = _898 & _912;
    assign _916 = write_enable_36 | read_enable_29;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_17
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_916), .regcea(vdd), .wea(write_enable_36), .addra(address_36), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_35), .regceb(vdd), .web(write_enable_35), .addrb(address_35), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_921[131:131]), .sbiterrb(_921[130:130]), .doutb(_921[129:66]), .dbiterra(_921[65:65]), .sbiterra(_921[64:64]), .douta(_921[63:0]) );
    assign _922 = _921[63:0];
    assign address_37 = PHASE_10 ? _199 : _907;
    assign _905 = _129 & _868;
    assign write_enable_37 = _905 & PHASE_10;
    assign _830 = _822[129:66];
    assign _829 = _809[129:66];
    assign _831 = PHASE_8 ? _830 : _829;
    assign _827 = _779[129:66];
    assign _826 = _765[129:66];
    assign q1_2 = PHASE_9 ? _827 : _826;
    assign _832 = _746 ? _831 : q1_2;
    assign address_38 = _811 ? _805 : _804;
    assign _817 = ~ _811;
    assign read_enable_30 = _102 & _817;
    assign address_39 = _811 ? _60 : _793;
    assign _813 = ~ _811;
    assign read_enable_31 = _102 & _813;
    assign _811 = ~ PHASE_8;
    assign write_enable_39 = _782 & _811;
    assign _815 = write_enable_39 | read_enable_31;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_18
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_815), .regcea(vdd), .wea(write_enable_39), .addra(address_39), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_30), .regceb(vdd), .web(write_enable_38), .addrb(address_38), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_822[131:131]), .sbiterrb(_822[130:130]), .doutb(_822[129:66]), .dbiterra(_822[65:65]), .sbiterra(_822[64:64]), .douta(_822[63:0]) );
    assign _823 = _822[63:0];
    assign _803 = _172[5:5];
    assign _802 = _172[4:4];
    assign _801 = _172[3:3];
    assign _800 = _172[2:2];
    assign _799 = _172[1:1];
    assign _798 = _172[0:0];
    assign _804 = { _798, _799, _800, _801, _802, _803 };
    assign address_40 = PHASE_8 ? _805 : _804;
    assign _795 = ~ PHASE_8;
    assign read_enable_32 = _102 & _795;
    assign data_37 = wr_d4;
    assign _792 = _137[5:5];
    assign _791 = _137[4:4];
    assign _790 = _137[3:3];
    assign _789 = _137[2:2];
    assign _788 = _137[1:1];
    assign _787 = _137[0:0];
    assign _793 = { _787, _788, _789, _790, _791, _792 };
    assign address_41 = PHASE_8 ? _60 : _793;
    assign _784 = ~ PHASE_8;
    assign read_enable_33 = _102 & _784;
    assign _782 = _62[4:4];
    assign write_enable_41 = _782 & PHASE_8;
    assign _786 = write_enable_41 | read_enable_33;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_19
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_786), .regcea(vdd), .wea(write_enable_41), .addra(address_41), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_32), .regceb(vdd), .web(write_enable_40), .addrb(address_40), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_809[131:131]), .sbiterrb(_809[130:130]), .doutb(_809[129:66]), .dbiterra(_809[65:65]), .sbiterra(_809[64:64]), .douta(_809[63:0]) );
    assign _810 = _809[63:0];
    assign _743 = ~ PHASE_8;
    assign _27 = _743;
    always @(posedge _84) begin
        if (_82)
            PHASE_8 <= _741;
        else
            if (_72)
                PHASE_8 <= _27;
    end
    assign _824 = PHASE_8 ? _823 : _810;
    assign address_42 = _767 ? _199 : _172;
    assign _774 = ~ _767;
    assign read_enable_34 = _102 & _774;
    assign write_enable_42 = _758 & _767;
    assign _776 = write_enable_42 | read_enable_34;
    assign address_43 = _767 ? _164 : _137;
    assign _769 = ~ _767;
    assign read_enable_35 = _102 & _769;
    assign _767 = ~ PHASE_9;
    assign write_enable_43 = _751 & _767;
    assign _771 = write_enable_43 | read_enable_35;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_20
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_771), .regcea(vdd), .wea(write_enable_43), .addra(address_43), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_776), .regceb(vdd), .web(write_enable_42), .addrb(address_42), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_779[131:131]), .sbiterrb(_779[130:130]), .doutb(_779[129:66]), .dbiterra(_779[65:65]), .sbiterra(_779[64:64]), .douta(_779[63:0]) );
    assign _780 = _779[63:0];
    assign _835 = _834[127:64];
    assign data_39 = _835;
    assign address_44 = PHASE_9 ? _199 : _172;
    assign _760 = ~ PHASE_9;
    assign read_enable_36 = _102 & _760;
    assign _757 = ~ _130;
    assign _758 = _129 & _757;
    assign write_enable_44 = _758 & PHASE_9;
    assign _762 = write_enable_44 | read_enable_36;
    assign address_45 = PHASE_9 ? _164 : _137;
    assign _753 = ~ PHASE_9;
    assign read_enable_37 = _102 & _753;
    assign _750 = ~ _130;
    assign _751 = _129 & _750;
    assign write_enable_45 = _751 & PHASE_9;
    assign _755 = write_enable_45 | read_enable_37;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_21
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_755), .regcea(vdd), .wea(write_enable_45), .addra(address_45), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_762), .regceb(vdd), .web(write_enable_44), .addrb(address_44), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_765[131:131]), .sbiterrb(_765[130:130]), .doutb(_765[129:66]), .dbiterra(_765[65:65]), .sbiterra(_765[64:64]), .douta(_765[63:0]) );
    assign _766 = _765[63:0];
    assign _836 = ~ PHASE_9;
    assign _29 = _836;
    always @(posedge _84) begin
        if (_82)
            PHASE_9 <= _748;
        else
            if (_99)
                PHASE_9 <= _29;
    end
    assign q0_2 = PHASE_9 ? _780 : _766;
    always @(posedge _84) begin
        if (_82)
            _746 <= _745;
        else
            _746 <= _92;
    end
    assign _825 = _746 ? _824 : q0_2;
    dp_19
        dp_3
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_825), .d2(_832), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_834[191:128]), .q2(_834[127:64]), .q1(_834[63:0]) );
    assign _837 = _834[63:0];
    assign data_43 = _837;
    assign address_46 = PHASE_10 ? _164 : _68;
    assign _901 = ~ PHASE_10;
    assign _900 = _70[4:4];
    assign read_enable_38 = _900 & _901;
    always @(posedge _84) begin
        if (_82)
            _871 <= _870;
        else
            _871 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _874 <= _873;
        else
            _874 <= _871;
    end
    always @(posedge _84) begin
        if (_82)
            _877 <= _876;
        else
            _877 <= _874;
    end
    always @(posedge _84) begin
        if (_82)
            _880 <= _879;
        else
            _880 <= _877;
    end
    always @(posedge _84) begin
        if (_82)
            _883 <= _882;
        else
            _883 <= _880;
    end
    always @(posedge _84) begin
        if (_82)
            _886 <= _885;
        else
            _886 <= _883;
    end
    always @(posedge _84) begin
        if (_82)
            _889 <= _888;
        else
            _889 <= _886;
    end
    always @(posedge _84) begin
        if (_82)
            _892 <= _891;
        else
            _892 <= _889;
    end
    always @(posedge _84) begin
        if (_82)
            _895 <= _894;
        else
            _895 <= _892;
    end
    assign _896 = ~ _895;
    always @(posedge _84) begin
        if (_82)
            _844 <= _843;
        else
            _844 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _847 <= _846;
        else
            _847 <= _844;
    end
    always @(posedge _84) begin
        if (_82)
            _850 <= _849;
        else
            _850 <= _847;
    end
    always @(posedge _84) begin
        if (_82)
            _853 <= _852;
        else
            _853 <= _850;
    end
    always @(posedge _84) begin
        if (_82)
            _856 <= _855;
        else
            _856 <= _853;
    end
    always @(posedge _84) begin
        if (_82)
            _859 <= _858;
        else
            _859 <= _856;
    end
    always @(posedge _84) begin
        if (_82)
            _862 <= _861;
        else
            _862 <= _859;
    end
    always @(posedge _84) begin
        if (_82)
            _865 <= _864;
        else
            _865 <= _862;
    end
    always @(posedge _84) begin
        if (_82)
            _868 <= _867;
        else
            _868 <= _865;
    end
    assign _897 = _868 & _896;
    assign _898 = _129 & _897;
    assign write_enable_46 = _898 & PHASE_10;
    assign _903 = write_enable_46 | read_enable_38;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_22
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_903), .regcea(vdd), .wea(write_enable_46), .addra(address_46), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_37), .regceb(vdd), .web(write_enable_37), .addrb(address_37), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_910[131:131]), .sbiterrb(_910[130:130]), .doutb(_910[129:66]), .dbiterra(_910[65:65]), .sbiterra(_910[64:64]), .douta(_910[63:0]) );
    assign _911 = _910[63:0];
    assign _841 = ~ PHASE_10;
    assign _31 = _841;
    always @(posedge _84) begin
        if (_82)
            PHASE_10 <= _839;
        else
            if (_72)
                PHASE_10 <= _31;
    end
    assign _923 = PHASE_10 ? _922 : _911;
    assign address_47 = _1096 ? _199 : _1091;
    assign write_enable_47 = _1089 & _1096;
    assign address_48 = _1096 ? _164 : _68;
    assign _1098 = ~ _1096;
    assign read_enable_39 = _1084 & _1098;
    assign _1096 = ~ PHASE_13;
    assign write_enable_48 = _1082 & _1096;
    assign _1100 = write_enable_48 | read_enable_39;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_23
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1100), .regcea(vdd), .wea(write_enable_48), .addra(address_48), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_47), .regceb(vdd), .web(write_enable_47), .addrb(address_47), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1105[131:131]), .sbiterrb(_1105[130:130]), .doutb(_1105[129:66]), .dbiterra(_1105[65:65]), .sbiterra(_1105[64:64]), .douta(_1105[63:0]) );
    assign _1106 = _1105[63:0];
    assign address_49 = PHASE_13 ? _199 : _1091;
    assign _1089 = _129 & _1052;
    assign write_enable_49 = _1089 & PHASE_13;
    assign _1014 = _1006[129:66];
    assign _1013 = _993[129:66];
    assign _1015 = PHASE_11 ? _1014 : _1013;
    assign _1011 = _963[129:66];
    assign _1010 = _949[129:66];
    assign q1_3 = PHASE_12 ? _1011 : _1010;
    assign _1016 = _930 ? _1015 : q1_3;
    assign address_50 = _995 ? _989 : _988;
    assign _1001 = ~ _995;
    assign read_enable_40 = _102 & _1001;
    assign address_51 = _995 ? _60 : _977;
    assign _997 = ~ _995;
    assign read_enable_41 = _102 & _997;
    assign _995 = ~ PHASE_11;
    assign write_enable_51 = _966 & _995;
    assign _999 = write_enable_51 | read_enable_41;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_24
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_999), .regcea(vdd), .wea(write_enable_51), .addra(address_51), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_40), .regceb(vdd), .web(write_enable_50), .addrb(address_50), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1006[131:131]), .sbiterrb(_1006[130:130]), .doutb(_1006[129:66]), .dbiterra(_1006[65:65]), .sbiterra(_1006[64:64]), .douta(_1006[63:0]) );
    assign _1007 = _1006[63:0];
    assign _987 = _172[5:5];
    assign _986 = _172[4:4];
    assign _985 = _172[3:3];
    assign _984 = _172[2:2];
    assign _983 = _172[1:1];
    assign _982 = _172[0:0];
    assign _988 = { _982, _983, _984, _985, _986, _987 };
    assign address_52 = PHASE_11 ? _989 : _988;
    assign _979 = ~ PHASE_11;
    assign read_enable_42 = _102 & _979;
    assign data_49 = wr_d3;
    assign _976 = _137[5:5];
    assign _975 = _137[4:4];
    assign _974 = _137[3:3];
    assign _973 = _137[2:2];
    assign _972 = _137[1:1];
    assign _971 = _137[0:0];
    assign _977 = { _971, _972, _973, _974, _975, _976 };
    assign address_53 = PHASE_11 ? _60 : _977;
    assign _968 = ~ PHASE_11;
    assign read_enable_43 = _102 & _968;
    assign _966 = _62[3:3];
    assign write_enable_53 = _966 & PHASE_11;
    assign _970 = write_enable_53 | read_enable_43;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_25
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_970), .regcea(vdd), .wea(write_enable_53), .addra(address_53), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_42), .regceb(vdd), .web(write_enable_52), .addrb(address_52), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_993[131:131]), .sbiterrb(_993[130:130]), .doutb(_993[129:66]), .dbiterra(_993[65:65]), .sbiterra(_993[64:64]), .douta(_993[63:0]) );
    assign _994 = _993[63:0];
    assign _927 = ~ PHASE_11;
    assign _35 = _927;
    always @(posedge _84) begin
        if (_82)
            PHASE_11 <= _925;
        else
            if (_72)
                PHASE_11 <= _35;
    end
    assign _1008 = PHASE_11 ? _1007 : _994;
    assign address_54 = _951 ? _199 : _172;
    assign _958 = ~ _951;
    assign read_enable_44 = _102 & _958;
    assign write_enable_54 = _942 & _951;
    assign _960 = write_enable_54 | read_enable_44;
    assign address_55 = _951 ? _164 : _137;
    assign _953 = ~ _951;
    assign read_enable_45 = _102 & _953;
    assign _951 = ~ PHASE_12;
    assign write_enable_55 = _935 & _951;
    assign _955 = write_enable_55 | read_enable_45;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_26
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_955), .regcea(vdd), .wea(write_enable_55), .addra(address_55), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_960), .regceb(vdd), .web(write_enable_54), .addrb(address_54), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_963[131:131]), .sbiterrb(_963[130:130]), .doutb(_963[129:66]), .dbiterra(_963[65:65]), .sbiterra(_963[64:64]), .douta(_963[63:0]) );
    assign _964 = _963[63:0];
    assign _1019 = _1018[127:64];
    assign data_51 = _1019;
    assign address_56 = PHASE_12 ? _199 : _172;
    assign _944 = ~ PHASE_12;
    assign read_enable_46 = _102 & _944;
    assign _941 = ~ _130;
    assign _942 = _129 & _941;
    assign write_enable_56 = _942 & PHASE_12;
    assign _946 = write_enable_56 | read_enable_46;
    assign address_57 = PHASE_12 ? _164 : _137;
    assign _937 = ~ PHASE_12;
    assign read_enable_47 = _102 & _937;
    assign _934 = ~ _130;
    assign _935 = _129 & _934;
    assign write_enable_57 = _935 & PHASE_12;
    assign _939 = write_enable_57 | read_enable_47;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_27
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_939), .regcea(vdd), .wea(write_enable_57), .addra(address_57), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_946), .regceb(vdd), .web(write_enable_56), .addrb(address_56), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_949[131:131]), .sbiterrb(_949[130:130]), .doutb(_949[129:66]), .dbiterra(_949[65:65]), .sbiterra(_949[64:64]), .douta(_949[63:0]) );
    assign _950 = _949[63:0];
    assign _1020 = ~ PHASE_12;
    assign _37 = _1020;
    always @(posedge _84) begin
        if (_82)
            PHASE_12 <= _932;
        else
            if (_99)
                PHASE_12 <= _37;
    end
    assign q0_3 = PHASE_12 ? _964 : _950;
    always @(posedge _84) begin
        if (_82)
            _930 <= _929;
        else
            _930 <= _92;
    end
    assign _1009 = _930 ? _1008 : q0_3;
    dp_18
        dp_2
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1009), .d2(_1016), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_1018[191:128]), .q2(_1018[127:64]), .q1(_1018[63:0]) );
    assign _1021 = _1018[63:0];
    assign data_55 = _1021;
    assign address_58 = PHASE_13 ? _164 : _68;
    assign _1085 = ~ PHASE_13;
    assign _1084 = _70[3:3];
    assign read_enable_48 = _1084 & _1085;
    always @(posedge _84) begin
        if (_82)
            _1055 <= _1054;
        else
            _1055 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _1058 <= _1057;
        else
            _1058 <= _1055;
    end
    always @(posedge _84) begin
        if (_82)
            _1061 <= _1060;
        else
            _1061 <= _1058;
    end
    always @(posedge _84) begin
        if (_82)
            _1064 <= _1063;
        else
            _1064 <= _1061;
    end
    always @(posedge _84) begin
        if (_82)
            _1067 <= _1066;
        else
            _1067 <= _1064;
    end
    always @(posedge _84) begin
        if (_82)
            _1070 <= _1069;
        else
            _1070 <= _1067;
    end
    always @(posedge _84) begin
        if (_82)
            _1073 <= _1072;
        else
            _1073 <= _1070;
    end
    always @(posedge _84) begin
        if (_82)
            _1076 <= _1075;
        else
            _1076 <= _1073;
    end
    always @(posedge _84) begin
        if (_82)
            _1079 <= _1078;
        else
            _1079 <= _1076;
    end
    assign _1080 = ~ _1079;
    always @(posedge _84) begin
        if (_82)
            _1028 <= _1027;
        else
            _1028 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1031 <= _1030;
        else
            _1031 <= _1028;
    end
    always @(posedge _84) begin
        if (_82)
            _1034 <= _1033;
        else
            _1034 <= _1031;
    end
    always @(posedge _84) begin
        if (_82)
            _1037 <= _1036;
        else
            _1037 <= _1034;
    end
    always @(posedge _84) begin
        if (_82)
            _1040 <= _1039;
        else
            _1040 <= _1037;
    end
    always @(posedge _84) begin
        if (_82)
            _1043 <= _1042;
        else
            _1043 <= _1040;
    end
    always @(posedge _84) begin
        if (_82)
            _1046 <= _1045;
        else
            _1046 <= _1043;
    end
    always @(posedge _84) begin
        if (_82)
            _1049 <= _1048;
        else
            _1049 <= _1046;
    end
    always @(posedge _84) begin
        if (_82)
            _1052 <= _1051;
        else
            _1052 <= _1049;
    end
    assign _1081 = _1052 & _1080;
    assign _1082 = _129 & _1081;
    assign write_enable_58 = _1082 & PHASE_13;
    assign _1087 = write_enable_58 | read_enable_48;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_28
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1087), .regcea(vdd), .wea(write_enable_58), .addra(address_58), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_49), .regceb(vdd), .web(write_enable_49), .addrb(address_49), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1094[131:131]), .sbiterrb(_1094[130:130]), .doutb(_1094[129:66]), .dbiterra(_1094[65:65]), .sbiterra(_1094[64:64]), .douta(_1094[63:0]) );
    assign _1095 = _1094[63:0];
    assign _1025 = ~ PHASE_13;
    assign _39 = _1025;
    always @(posedge _84) begin
        if (_82)
            PHASE_13 <= _1023;
        else
            if (_72)
                PHASE_13 <= _39;
    end
    assign _1107 = PHASE_13 ? _1106 : _1095;
    assign address_59 = _1280 ? _199 : _1275;
    assign write_enable_59 = _1273 & _1280;
    assign address_60 = _1280 ? _164 : _68;
    assign _1282 = ~ _1280;
    assign read_enable_49 = _1268 & _1282;
    assign _1280 = ~ PHASE_16;
    assign write_enable_60 = _1266 & _1280;
    assign _1284 = write_enable_60 | read_enable_49;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_29
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1284), .regcea(vdd), .wea(write_enable_60), .addra(address_60), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_59), .regceb(vdd), .web(write_enable_59), .addrb(address_59), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1289[131:131]), .sbiterrb(_1289[130:130]), .doutb(_1289[129:66]), .dbiterra(_1289[65:65]), .sbiterra(_1289[64:64]), .douta(_1289[63:0]) );
    assign _1290 = _1289[63:0];
    assign address_61 = PHASE_16 ? _199 : _1275;
    assign _1273 = _129 & _1236;
    assign write_enable_61 = _1273 & PHASE_16;
    assign _1198 = _1190[129:66];
    assign _1197 = _1177[129:66];
    assign _1199 = PHASE_14 ? _1198 : _1197;
    assign _1195 = _1147[129:66];
    assign _1194 = _1133[129:66];
    assign q1_4 = PHASE_15 ? _1195 : _1194;
    assign _1200 = _1114 ? _1199 : q1_4;
    assign address_62 = _1179 ? _1173 : _1172;
    assign _1185 = ~ _1179;
    assign read_enable_50 = _102 & _1185;
    assign address_63 = _1179 ? _60 : _1161;
    assign _1181 = ~ _1179;
    assign read_enable_51 = _102 & _1181;
    assign _1179 = ~ PHASE_14;
    assign write_enable_63 = _1150 & _1179;
    assign _1183 = write_enable_63 | read_enable_51;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_30
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1183), .regcea(vdd), .wea(write_enable_63), .addra(address_63), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_50), .regceb(vdd), .web(write_enable_62), .addrb(address_62), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1190[131:131]), .sbiterrb(_1190[130:130]), .doutb(_1190[129:66]), .dbiterra(_1190[65:65]), .sbiterra(_1190[64:64]), .douta(_1190[63:0]) );
    assign _1191 = _1190[63:0];
    assign _1171 = _172[5:5];
    assign _1170 = _172[4:4];
    assign _1169 = _172[3:3];
    assign _1168 = _172[2:2];
    assign _1167 = _172[1:1];
    assign _1166 = _172[0:0];
    assign _1172 = { _1166, _1167, _1168, _1169, _1170, _1171 };
    assign address_64 = PHASE_14 ? _1173 : _1172;
    assign _1163 = ~ PHASE_14;
    assign read_enable_52 = _102 & _1163;
    assign data_61 = wr_d2;
    assign _1160 = _137[5:5];
    assign _1159 = _137[4:4];
    assign _1158 = _137[3:3];
    assign _1157 = _137[2:2];
    assign _1156 = _137[1:1];
    assign _1155 = _137[0:0];
    assign _1161 = { _1155, _1156, _1157, _1158, _1159, _1160 };
    assign address_65 = PHASE_14 ? _60 : _1161;
    assign _1152 = ~ PHASE_14;
    assign read_enable_53 = _102 & _1152;
    assign _1150 = _62[2:2];
    assign write_enable_65 = _1150 & PHASE_14;
    assign _1154 = write_enable_65 | read_enable_53;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_31
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1154), .regcea(vdd), .wea(write_enable_65), .addra(address_65), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_52), .regceb(vdd), .web(write_enable_64), .addrb(address_64), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1177[131:131]), .sbiterrb(_1177[130:130]), .doutb(_1177[129:66]), .dbiterra(_1177[65:65]), .sbiterra(_1177[64:64]), .douta(_1177[63:0]) );
    assign _1178 = _1177[63:0];
    assign _1111 = ~ PHASE_14;
    assign _43 = _1111;
    always @(posedge _84) begin
        if (_82)
            PHASE_14 <= _1109;
        else
            if (_72)
                PHASE_14 <= _43;
    end
    assign _1192 = PHASE_14 ? _1191 : _1178;
    assign address_66 = _1135 ? _199 : _172;
    assign _1142 = ~ _1135;
    assign read_enable_54 = _102 & _1142;
    assign write_enable_66 = _1126 & _1135;
    assign _1144 = write_enable_66 | read_enable_54;
    assign address_67 = _1135 ? _164 : _137;
    assign _1137 = ~ _1135;
    assign read_enable_55 = _102 & _1137;
    assign _1135 = ~ PHASE_15;
    assign write_enable_67 = _1119 & _1135;
    assign _1139 = write_enable_67 | read_enable_55;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_32
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1139), .regcea(vdd), .wea(write_enable_67), .addra(address_67), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1144), .regceb(vdd), .web(write_enable_66), .addrb(address_66), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1147[131:131]), .sbiterrb(_1147[130:130]), .doutb(_1147[129:66]), .dbiterra(_1147[65:65]), .sbiterra(_1147[64:64]), .douta(_1147[63:0]) );
    assign _1148 = _1147[63:0];
    assign _1203 = _1202[127:64];
    assign data_63 = _1203;
    assign address_68 = PHASE_15 ? _199 : _172;
    assign _1128 = ~ PHASE_15;
    assign read_enable_56 = _102 & _1128;
    assign _1125 = ~ _130;
    assign _1126 = _129 & _1125;
    assign write_enable_68 = _1126 & PHASE_15;
    assign _1130 = write_enable_68 | read_enable_56;
    assign address_69 = PHASE_15 ? _164 : _137;
    assign _1121 = ~ PHASE_15;
    assign read_enable_57 = _102 & _1121;
    assign _1118 = ~ _130;
    assign _1119 = _129 & _1118;
    assign write_enable_69 = _1119 & PHASE_15;
    assign _1123 = write_enable_69 | read_enable_57;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_33
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1123), .regcea(vdd), .wea(write_enable_69), .addra(address_69), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1130), .regceb(vdd), .web(write_enable_68), .addrb(address_68), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1133[131:131]), .sbiterrb(_1133[130:130]), .doutb(_1133[129:66]), .dbiterra(_1133[65:65]), .sbiterra(_1133[64:64]), .douta(_1133[63:0]) );
    assign _1134 = _1133[63:0];
    assign _1204 = ~ PHASE_15;
    assign _45 = _1204;
    always @(posedge _84) begin
        if (_82)
            PHASE_15 <= _1116;
        else
            if (_99)
                PHASE_15 <= _45;
    end
    assign q0_4 = PHASE_15 ? _1148 : _1134;
    always @(posedge _84) begin
        if (_82)
            _1114 <= _1113;
        else
            _1114 <= _92;
    end
    assign _1193 = _1114 ? _1192 : q0_4;
    dp_17
        dp_1
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1193), .d2(_1200), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_1202[191:128]), .q2(_1202[127:64]), .q1(_1202[63:0]) );
    assign _1205 = _1202[63:0];
    assign data_67 = _1205;
    assign address_70 = PHASE_16 ? _164 : _68;
    assign _1269 = ~ PHASE_16;
    assign _1268 = _70[2:2];
    assign read_enable_58 = _1268 & _1269;
    always @(posedge _84) begin
        if (_82)
            _1239 <= _1238;
        else
            _1239 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _1242 <= _1241;
        else
            _1242 <= _1239;
    end
    always @(posedge _84) begin
        if (_82)
            _1245 <= _1244;
        else
            _1245 <= _1242;
    end
    always @(posedge _84) begin
        if (_82)
            _1248 <= _1247;
        else
            _1248 <= _1245;
    end
    always @(posedge _84) begin
        if (_82)
            _1251 <= _1250;
        else
            _1251 <= _1248;
    end
    always @(posedge _84) begin
        if (_82)
            _1254 <= _1253;
        else
            _1254 <= _1251;
    end
    always @(posedge _84) begin
        if (_82)
            _1257 <= _1256;
        else
            _1257 <= _1254;
    end
    always @(posedge _84) begin
        if (_82)
            _1260 <= _1259;
        else
            _1260 <= _1257;
    end
    always @(posedge _84) begin
        if (_82)
            _1263 <= _1262;
        else
            _1263 <= _1260;
    end
    assign _1264 = ~ _1263;
    always @(posedge _84) begin
        if (_82)
            _1212 <= _1211;
        else
            _1212 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1215 <= _1214;
        else
            _1215 <= _1212;
    end
    always @(posedge _84) begin
        if (_82)
            _1218 <= _1217;
        else
            _1218 <= _1215;
    end
    always @(posedge _84) begin
        if (_82)
            _1221 <= _1220;
        else
            _1221 <= _1218;
    end
    always @(posedge _84) begin
        if (_82)
            _1224 <= _1223;
        else
            _1224 <= _1221;
    end
    always @(posedge _84) begin
        if (_82)
            _1227 <= _1226;
        else
            _1227 <= _1224;
    end
    always @(posedge _84) begin
        if (_82)
            _1230 <= _1229;
        else
            _1230 <= _1227;
    end
    always @(posedge _84) begin
        if (_82)
            _1233 <= _1232;
        else
            _1233 <= _1230;
    end
    always @(posedge _84) begin
        if (_82)
            _1236 <= _1235;
        else
            _1236 <= _1233;
    end
    assign _1265 = _1236 & _1264;
    assign _1266 = _129 & _1265;
    assign write_enable_70 = _1266 & PHASE_16;
    assign _1271 = write_enable_70 | read_enable_58;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_34
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1271), .regcea(vdd), .wea(write_enable_70), .addra(address_70), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_61), .regceb(vdd), .web(write_enable_61), .addrb(address_61), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1278[131:131]), .sbiterrb(_1278[130:130]), .doutb(_1278[129:66]), .dbiterra(_1278[65:65]), .sbiterra(_1278[64:64]), .douta(_1278[63:0]) );
    assign _1279 = _1278[63:0];
    assign _1209 = ~ PHASE_16;
    assign _47 = _1209;
    always @(posedge _84) begin
        if (_82)
            PHASE_16 <= _1207;
        else
            if (_72)
                PHASE_16 <= _47;
    end
    assign _1291 = PHASE_16 ? _1290 : _1279;
    assign address_71 = _1464 ? _199 : _1459;
    assign write_enable_71 = _1457 & _1464;
    assign address_72 = _1464 ? _164 : _68;
    assign _1466 = ~ _1464;
    assign read_enable_59 = _1452 & _1466;
    assign _1464 = ~ PHASE_19;
    assign write_enable_72 = _1450 & _1464;
    assign _1468 = write_enable_72 | read_enable_59;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_35
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1468), .regcea(vdd), .wea(write_enable_72), .addra(address_72), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_71), .regceb(vdd), .web(write_enable_71), .addrb(address_71), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1473[131:131]), .sbiterrb(_1473[130:130]), .doutb(_1473[129:66]), .dbiterra(_1473[65:65]), .sbiterra(_1473[64:64]), .douta(_1473[63:0]) );
    assign _1474 = _1473[63:0];
    assign address_73 = PHASE_19 ? _199 : _1459;
    assign _1457 = _129 & _1420;
    assign write_enable_73 = _1457 & PHASE_19;
    assign _1382 = _1374[129:66];
    assign _1381 = _1361[129:66];
    assign _1383 = PHASE_17 ? _1382 : _1381;
    assign _1379 = _1331[129:66];
    assign _1378 = _1317[129:66];
    assign q1_5 = PHASE_18 ? _1379 : _1378;
    assign _1384 = _1298 ? _1383 : q1_5;
    assign address_74 = _1363 ? _1357 : _1356;
    assign _1369 = ~ _1363;
    assign read_enable_60 = _102 & _1369;
    assign address_75 = _1363 ? _60 : _1345;
    assign _1365 = ~ _1363;
    assign read_enable_61 = _102 & _1365;
    assign _1363 = ~ PHASE_17;
    assign write_enable_75 = _1334 & _1363;
    assign _1367 = write_enable_75 | read_enable_61;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_36
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1367), .regcea(vdd), .wea(write_enable_75), .addra(address_75), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_60), .regceb(vdd), .web(write_enable_74), .addrb(address_74), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1374[131:131]), .sbiterrb(_1374[130:130]), .doutb(_1374[129:66]), .dbiterra(_1374[65:65]), .sbiterra(_1374[64:64]), .douta(_1374[63:0]) );
    assign _1375 = _1374[63:0];
    assign _1355 = _172[5:5];
    assign _1354 = _172[4:4];
    assign _1353 = _172[3:3];
    assign _1352 = _172[2:2];
    assign _1351 = _172[1:1];
    assign _1350 = _172[0:0];
    assign _1356 = { _1350, _1351, _1352, _1353, _1354, _1355 };
    assign address_76 = PHASE_17 ? _1357 : _1356;
    assign _1347 = ~ PHASE_17;
    assign read_enable_62 = _102 & _1347;
    assign data_73 = wr_d1;
    assign _1344 = _137[5:5];
    assign _1343 = _137[4:4];
    assign _1342 = _137[3:3];
    assign _1341 = _137[2:2];
    assign _1340 = _137[1:1];
    assign _1339 = _137[0:0];
    assign _1345 = { _1339, _1340, _1341, _1342, _1343, _1344 };
    assign address_77 = PHASE_17 ? _60 : _1345;
    assign _1336 = ~ PHASE_17;
    assign read_enable_63 = _102 & _1336;
    assign _1334 = _62[1:1];
    assign write_enable_77 = _1334 & PHASE_17;
    assign _1338 = write_enable_77 | read_enable_63;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_37
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1338), .regcea(vdd), .wea(write_enable_77), .addra(address_77), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_62), .regceb(vdd), .web(write_enable_76), .addrb(address_76), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1361[131:131]), .sbiterrb(_1361[130:130]), .doutb(_1361[129:66]), .dbiterra(_1361[65:65]), .sbiterra(_1361[64:64]), .douta(_1361[63:0]) );
    assign _1362 = _1361[63:0];
    assign _1295 = ~ PHASE_17;
    assign _51 = _1295;
    always @(posedge _84) begin
        if (_82)
            PHASE_17 <= _1293;
        else
            if (_72)
                PHASE_17 <= _51;
    end
    assign _1376 = PHASE_17 ? _1375 : _1362;
    assign address_78 = _1319 ? _199 : _172;
    assign _1326 = ~ _1319;
    assign read_enable_64 = _102 & _1326;
    assign write_enable_78 = _1310 & _1319;
    assign _1328 = write_enable_78 | read_enable_64;
    assign address_79 = _1319 ? _164 : _137;
    assign _1321 = ~ _1319;
    assign read_enable_65 = _102 & _1321;
    assign _1319 = ~ PHASE_18;
    assign write_enable_79 = _1303 & _1319;
    assign _1323 = write_enable_79 | read_enable_65;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_38
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1323), .regcea(vdd), .wea(write_enable_79), .addra(address_79), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1328), .regceb(vdd), .web(write_enable_78), .addrb(address_78), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1331[131:131]), .sbiterrb(_1331[130:130]), .doutb(_1331[129:66]), .dbiterra(_1331[65:65]), .sbiterra(_1331[64:64]), .douta(_1331[63:0]) );
    assign _1332 = _1331[63:0];
    assign _1387 = _1386[127:64];
    assign data_75 = _1387;
    assign address_80 = PHASE_18 ? _199 : _172;
    assign _1312 = ~ PHASE_18;
    assign read_enable_66 = _102 & _1312;
    assign _1309 = ~ _130;
    assign _1310 = _129 & _1309;
    assign write_enable_80 = _1310 & PHASE_18;
    assign _1314 = write_enable_80 | read_enable_66;
    assign address_81 = PHASE_18 ? _164 : _137;
    assign _1305 = ~ PHASE_18;
    assign read_enable_67 = _102 & _1305;
    assign _1302 = ~ _130;
    assign _1303 = _129 & _1302;
    assign write_enable_81 = _1303 & PHASE_18;
    assign _1307 = write_enable_81 | read_enable_67;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_39
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1307), .regcea(vdd), .wea(write_enable_81), .addra(address_81), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1314), .regceb(vdd), .web(write_enable_80), .addrb(address_80), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1317[131:131]), .sbiterrb(_1317[130:130]), .doutb(_1317[129:66]), .dbiterra(_1317[65:65]), .sbiterra(_1317[64:64]), .douta(_1317[63:0]) );
    assign _1318 = _1317[63:0];
    assign _1388 = ~ PHASE_18;
    assign _53 = _1388;
    always @(posedge _84) begin
        if (_82)
            PHASE_18 <= _1300;
        else
            if (_99)
                PHASE_18 <= _53;
    end
    assign q0_5 = PHASE_18 ? _1332 : _1318;
    always @(posedge _84) begin
        if (_82)
            _1298 <= _1297;
        else
            _1298 <= _92;
    end
    assign _1377 = _1298 ? _1376 : q0_5;
    dp_16
        dp_0
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1377), .d2(_1384), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_1386[191:128]), .q2(_1386[127:64]), .q1(_1386[63:0]) );
    assign _1389 = _1386[63:0];
    assign data_79 = _1389;
    assign address_82 = PHASE_19 ? _164 : _68;
    assign _1453 = ~ PHASE_19;
    assign _1452 = _70[1:1];
    assign read_enable_68 = _1452 & _1453;
    always @(posedge _84) begin
        if (_82)
            _1423 <= _1422;
        else
            _1423 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _1426 <= _1425;
        else
            _1426 <= _1423;
    end
    always @(posedge _84) begin
        if (_82)
            _1429 <= _1428;
        else
            _1429 <= _1426;
    end
    always @(posedge _84) begin
        if (_82)
            _1432 <= _1431;
        else
            _1432 <= _1429;
    end
    always @(posedge _84) begin
        if (_82)
            _1435 <= _1434;
        else
            _1435 <= _1432;
    end
    always @(posedge _84) begin
        if (_82)
            _1438 <= _1437;
        else
            _1438 <= _1435;
    end
    always @(posedge _84) begin
        if (_82)
            _1441 <= _1440;
        else
            _1441 <= _1438;
    end
    always @(posedge _84) begin
        if (_82)
            _1444 <= _1443;
        else
            _1444 <= _1441;
    end
    always @(posedge _84) begin
        if (_82)
            _1447 <= _1446;
        else
            _1447 <= _1444;
    end
    assign _1448 = ~ _1447;
    always @(posedge _84) begin
        if (_82)
            _1396 <= _1395;
        else
            _1396 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1399 <= _1398;
        else
            _1399 <= _1396;
    end
    always @(posedge _84) begin
        if (_82)
            _1402 <= _1401;
        else
            _1402 <= _1399;
    end
    always @(posedge _84) begin
        if (_82)
            _1405 <= _1404;
        else
            _1405 <= _1402;
    end
    always @(posedge _84) begin
        if (_82)
            _1408 <= _1407;
        else
            _1408 <= _1405;
    end
    always @(posedge _84) begin
        if (_82)
            _1411 <= _1410;
        else
            _1411 <= _1408;
    end
    always @(posedge _84) begin
        if (_82)
            _1414 <= _1413;
        else
            _1414 <= _1411;
    end
    always @(posedge _84) begin
        if (_82)
            _1417 <= _1416;
        else
            _1417 <= _1414;
    end
    always @(posedge _84) begin
        if (_82)
            _1420 <= _1419;
        else
            _1420 <= _1417;
    end
    assign _1449 = _1420 & _1448;
    assign _1450 = _129 & _1449;
    assign write_enable_82 = _1450 & PHASE_19;
    assign _1455 = write_enable_82 | read_enable_68;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_40
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1455), .regcea(vdd), .wea(write_enable_82), .addra(address_82), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_73), .regceb(vdd), .web(write_enable_73), .addrb(address_73), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1462[131:131]), .sbiterrb(_1462[130:130]), .doutb(_1462[129:66]), .dbiterra(_1462[65:65]), .sbiterra(_1462[64:64]), .douta(_1462[63:0]) );
    assign _1463 = _1462[63:0];
    assign _1393 = ~ PHASE_19;
    assign _55 = _1393;
    always @(posedge _84) begin
        if (_82)
            PHASE_19 <= _1391;
        else
            if (_72)
                PHASE_19 <= _55;
    end
    assign _1475 = PHASE_19 ? _1474 : _1463;
    assign address_83 = _1648 ? _199 : _1643;
    assign write_enable_83 = _1641 & _1648;
    assign address_84 = _1648 ? _164 : _68;
    assign _1650 = ~ _1648;
    assign read_enable_69 = _1636 & _1650;
    assign _1648 = ~ PHASE_22;
    assign write_enable_84 = _1634 & _1648;
    assign _1652 = write_enable_84 | read_enable_69;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_41
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1652), .regcea(vdd), .wea(write_enable_84), .addra(address_84), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_83), .regceb(vdd), .web(write_enable_83), .addrb(address_83), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1657[131:131]), .sbiterrb(_1657[130:130]), .doutb(_1657[129:66]), .dbiterra(_1657[65:65]), .sbiterra(_1657[64:64]), .douta(_1657[63:0]) );
    assign _1658 = _1657[63:0];
    assign address_85 = PHASE_22 ? _199 : _1643;
    assign _1641 = _129 & _1604;
    assign write_enable_85 = _1641 & PHASE_22;
    assign _280 = _91[490:487];
    assign _279 = _91[486:486];
    assign _277 = _91[482:482];
    assign _276 = _91[481:418];
    assign _275 = _91[417:354];
    assign _274 = _91[353:290];
    assign _273 = _91[289:226];
    assign _272 = _91[225:162];
    assign _271 = _91[161:98];
    assign _270 = _91[97:34];
    assign _1566 = _1558[129:66];
    assign _1565 = _1545[129:66];
    assign _1567 = PHASE_20 ? _1566 : _1565;
    assign _1563 = _1515[129:66];
    assign _1562 = _1501[129:66];
    assign q1_6 = PHASE_21 ? _1563 : _1562;
    assign _1568 = _1482 ? _1567 : q1_6;
    assign address_86 = _1547 ? _1541 : _1540;
    assign _1553 = ~ _1547;
    assign read_enable_70 = _102 & _1553;
    assign address_87 = _1547 ? _60 : _1529;
    assign _1549 = ~ _1547;
    assign read_enable_71 = _102 & _1549;
    assign _1547 = ~ PHASE_20;
    assign write_enable_87 = _1518 & _1547;
    assign _1551 = write_enable_87 | read_enable_71;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_42
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1551), .regcea(vdd), .wea(write_enable_87), .addra(address_87), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_70), .regceb(vdd), .web(write_enable_86), .addrb(address_86), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1558[131:131]), .sbiterrb(_1558[130:130]), .doutb(_1558[129:66]), .dbiterra(_1558[65:65]), .sbiterra(_1558[64:64]), .douta(_1558[63:0]) );
    assign _1559 = _1558[63:0];
    assign _1539 = _172[5:5];
    assign _1538 = _172[4:4];
    assign _1537 = _172[3:3];
    assign _1536 = _172[2:2];
    assign _1535 = _172[1:1];
    assign _1534 = _172[0:0];
    assign _1540 = { _1534, _1535, _1536, _1537, _1538, _1539 };
    assign address_88 = PHASE_20 ? _1541 : _1540;
    assign _1531 = ~ PHASE_20;
    assign read_enable_72 = _102 & _1531;
    assign data_85 = wr_d0;
    assign _60 = wr_addr;
    assign _1528 = _137[5:5];
    assign _1527 = _137[4:4];
    assign _1526 = _137[3:3];
    assign _1525 = _137[2:2];
    assign _1524 = _137[1:1];
    assign _1523 = _137[0:0];
    assign _1529 = { _1523, _1524, _1525, _1526, _1527, _1528 };
    assign address_89 = PHASE_20 ? _60 : _1529;
    assign _1520 = ~ PHASE_20;
    assign read_enable_73 = _102 & _1520;
    assign _62 = wr_en;
    assign _1518 = _62[0:0];
    assign write_enable_89 = _1518 & PHASE_20;
    assign _1522 = write_enable_89 | read_enable_73;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_43
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1522), .regcea(vdd), .wea(write_enable_89), .addra(address_89), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_72), .regceb(vdd), .web(write_enable_88), .addrb(address_88), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1545[131:131]), .sbiterrb(_1545[130:130]), .doutb(_1545[129:66]), .dbiterra(_1545[65:65]), .sbiterra(_1545[64:64]), .douta(_1545[63:0]) );
    assign _1546 = _1545[63:0];
    assign _1479 = ~ PHASE_20;
    assign _63 = _1479;
    always @(posedge _84) begin
        if (_82)
            PHASE_20 <= _1477;
        else
            if (_72)
                PHASE_20 <= _63;
    end
    assign _1560 = PHASE_20 ? _1559 : _1546;
    assign address_90 = _1503 ? _199 : _172;
    assign _1510 = ~ _1503;
    assign read_enable_74 = _102 & _1510;
    assign write_enable_90 = _1494 & _1503;
    assign _1512 = write_enable_90 | read_enable_74;
    assign address_91 = _1503 ? _164 : _137;
    assign _1505 = ~ _1503;
    assign read_enable_75 = _102 & _1505;
    assign _1503 = ~ PHASE_21;
    assign write_enable_91 = _1487 & _1503;
    assign _1507 = write_enable_91 | read_enable_75;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_44
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1507), .regcea(vdd), .wea(write_enable_91), .addra(address_91), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1512), .regceb(vdd), .web(write_enable_90), .addrb(address_90), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1515[131:131]), .sbiterrb(_1515[130:130]), .doutb(_1515[129:66]), .dbiterra(_1515[65:65]), .sbiterra(_1515[64:64]), .douta(_1515[63:0]) );
    assign _1516 = _1515[63:0];
    assign _1571 = _1570[127:64];
    assign data_87 = _1571;
    always @(posedge _84) begin
        if (_82)
            _175 <= _174;
        else
            _175 <= _172;
    end
    always @(posedge _84) begin
        if (_82)
            _178 <= _177;
        else
            _178 <= _175;
    end
    always @(posedge _84) begin
        if (_82)
            _181 <= _180;
        else
            _181 <= _178;
    end
    always @(posedge _84) begin
        if (_82)
            _184 <= _183;
        else
            _184 <= _181;
    end
    always @(posedge _84) begin
        if (_82)
            _187 <= _186;
        else
            _187 <= _184;
    end
    always @(posedge _84) begin
        if (_82)
            _190 <= _189;
        else
            _190 <= _187;
    end
    always @(posedge _84) begin
        if (_82)
            _193 <= _192;
        else
            _193 <= _190;
    end
    always @(posedge _84) begin
        if (_82)
            _196 <= _195;
        else
            _196 <= _193;
    end
    always @(posedge _84) begin
        if (_82)
            _199 <= _198;
        else
            _199 <= _196;
    end
    assign _172 = _91[33:28];
    assign address_92 = PHASE_21 ? _199 : _172;
    assign _1496 = ~ PHASE_21;
    assign read_enable_76 = _102 & _1496;
    assign _1493 = ~ _130;
    assign _1494 = _129 & _1493;
    assign write_enable_92 = _1494 & PHASE_21;
    assign _1498 = write_enable_92 | read_enable_76;
    assign address_93 = PHASE_21 ? _164 : _137;
    assign _1489 = ~ PHASE_21;
    assign read_enable_77 = _102 & _1489;
    assign _1486 = ~ _130;
    assign _1487 = _129 & _1486;
    assign write_enable_93 = _1487 & PHASE_21;
    assign _1491 = write_enable_93 | read_enable_77;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_45
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1491), .regcea(vdd), .wea(write_enable_93), .addra(address_93), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1498), .regceb(vdd), .web(write_enable_92), .addrb(address_92), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1501[131:131]), .sbiterrb(_1501[130:130]), .doutb(_1501[129:66]), .dbiterra(_1501[65:65]), .sbiterra(_1501[64:64]), .douta(_1501[63:0]) );
    assign _1502 = _1501[63:0];
    assign _99 = _91[492:492];
    assign _1572 = ~ PHASE_21;
    assign _65 = _1572;
    always @(posedge _84) begin
        if (_82)
            PHASE_21 <= _1484;
        else
            if (_99)
                PHASE_21 <= _65;
    end
    assign q0_6 = PHASE_21 ? _1516 : _1502;
    assign _92 = _91[483:483];
    always @(posedge _84) begin
        if (_82)
            _1482 <= _1481;
        else
            _1482 <= _92;
    end
    assign _1561 = _1482 ? _1560 : q0_6;
    dp_15
        dp
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1561), .d2(_1568), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_1570[191:128]), .q2(_1570[127:64]), .q1(_1570[63:0]) );
    assign _1573 = _1570[63:0];
    assign data_91 = _1573;
    assign _137 = _91[27:22];
    always @(posedge _84) begin
        if (_82)
            _140 <= _139;
        else
            _140 <= _137;
    end
    always @(posedge _84) begin
        if (_82)
            _143 <= _142;
        else
            _143 <= _140;
    end
    always @(posedge _84) begin
        if (_82)
            _146 <= _145;
        else
            _146 <= _143;
    end
    always @(posedge _84) begin
        if (_82)
            _149 <= _148;
        else
            _149 <= _146;
    end
    always @(posedge _84) begin
        if (_82)
            _152 <= _151;
        else
            _152 <= _149;
    end
    always @(posedge _84) begin
        if (_82)
            _155 <= _154;
        else
            _155 <= _152;
    end
    always @(posedge _84) begin
        if (_82)
            _158 <= _157;
        else
            _158 <= _155;
    end
    always @(posedge _84) begin
        if (_82)
            _161 <= _160;
        else
            _161 <= _158;
    end
    always @(posedge _84) begin
        if (_82)
            _164 <= _163;
        else
            _164 <= _161;
    end
    assign _68 = rd_addr;
    assign address_94 = PHASE_22 ? _164 : _68;
    assign _1637 = ~ PHASE_22;
    assign _70 = rd_en;
    assign _1636 = _70[0:0];
    assign read_enable_78 = _1636 & _1637;
    assign _278 = _91[485:485];
    always @(posedge _84) begin
        if (_82)
            _1607 <= _1606;
        else
            _1607 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _1610 <= _1609;
        else
            _1610 <= _1607;
    end
    always @(posedge _84) begin
        if (_82)
            _1613 <= _1612;
        else
            _1613 <= _1610;
    end
    always @(posedge _84) begin
        if (_82)
            _1616 <= _1615;
        else
            _1616 <= _1613;
    end
    always @(posedge _84) begin
        if (_82)
            _1619 <= _1618;
        else
            _1619 <= _1616;
    end
    always @(posedge _84) begin
        if (_82)
            _1622 <= _1621;
        else
            _1622 <= _1619;
    end
    always @(posedge _84) begin
        if (_82)
            _1625 <= _1624;
        else
            _1625 <= _1622;
    end
    always @(posedge _84) begin
        if (_82)
            _1628 <= _1627;
        else
            _1628 <= _1625;
    end
    always @(posedge _84) begin
        if (_82)
            _1631 <= _1630;
        else
            _1631 <= _1628;
    end
    assign _1632 = ~ _1631;
    assign _130 = _91[484:484];
    always @(posedge _84) begin
        if (_82)
            _1580 <= _1579;
        else
            _1580 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1583 <= _1582;
        else
            _1583 <= _1580;
    end
    always @(posedge _84) begin
        if (_82)
            _1586 <= _1585;
        else
            _1586 <= _1583;
    end
    always @(posedge _84) begin
        if (_82)
            _1589 <= _1588;
        else
            _1589 <= _1586;
    end
    always @(posedge _84) begin
        if (_82)
            _1592 <= _1591;
        else
            _1592 <= _1589;
    end
    always @(posedge _84) begin
        if (_82)
            _1595 <= _1594;
        else
            _1595 <= _1592;
    end
    always @(posedge _84) begin
        if (_82)
            _1598 <= _1597;
        else
            _1598 <= _1595;
    end
    always @(posedge _84) begin
        if (_82)
            _1601 <= _1600;
        else
            _1601 <= _1598;
    end
    always @(posedge _84) begin
        if (_82)
            _1604 <= _1603;
        else
            _1604 <= _1601;
    end
    assign _1633 = _1604 & _1632;
    assign _102 = _91[491:491];
    always @(posedge _84) begin
        if (_82)
            _105 <= _104;
        else
            _105 <= _102;
    end
    always @(posedge _84) begin
        if (_82)
            _108 <= _107;
        else
            _108 <= _105;
    end
    always @(posedge _84) begin
        if (_82)
            _111 <= _110;
        else
            _111 <= _108;
    end
    always @(posedge _84) begin
        if (_82)
            _114 <= _113;
        else
            _114 <= _111;
    end
    always @(posedge _84) begin
        if (_82)
            _117 <= _116;
        else
            _117 <= _114;
    end
    always @(posedge _84) begin
        if (_82)
            _120 <= _119;
        else
            _120 <= _117;
    end
    always @(posedge _84) begin
        if (_82)
            _123 <= _122;
        else
            _123 <= _120;
    end
    always @(posedge _84) begin
        if (_82)
            _126 <= _125;
        else
            _126 <= _123;
    end
    always @(posedge _84) begin
        if (_82)
            _129 <= _128;
        else
            _129 <= _126;
    end
    assign _1634 = _129 & _1633;
    assign write_enable_94 = _1634 & PHASE_22;
    assign _1639 = write_enable_94 | read_enable_78;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_46
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1639), .regcea(vdd), .wea(write_enable_94), .addra(address_94), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_85), .regceb(vdd), .web(write_enable_85), .addrb(address_85), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1646[131:131]), .sbiterrb(_1646[130:130]), .doutb(_1646[129:66]), .dbiterra(_1646[65:65]), .sbiterra(_1646[64:64]), .douta(_1646[63:0]) );
    assign _1647 = _1646[63:0];
    assign _72 = flip;
    assign _1577 = ~ PHASE_22;
    assign _73 = _1577;
    always @(posedge _84) begin
        if (_82)
            PHASE_22 <= _1575;
        else
            if (_72)
                PHASE_22 <= _73;
    end
    assign _1659 = PHASE_22 ? _1658 : _1647;
    assign _76 = first_4step_pass;
    assign _78 = first_iter;
    assign _80 = start;
    assign _82 = clear;
    assign _84 = clock;
    ctrl
        ctrl
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .first_4step_pass(_76), .flip(_91[492:492]), .read_write_enable(_91[491:491]), .index(_91[490:487]), .valid(_91[486:486]), .twiddle_stage(_91[485:485]), .last_stage(_91[484:484]), .first_stage(_91[483:483]), .start_twiddles(_91[482:482]), .omegas6(_91[481:418]), .omegas5(_91[417:354]), .omegas4(_91[353:290]), .omegas3(_91[289:226]), .omegas2(_91[225:162]), .omegas1(_91[161:98]), .omegas0(_91[97:34]), .addr2(_91[33:28]), .addr1(_91[27:22]), .m(_91[21:16]), .k(_91[15:10]), .j(_91[9:4]), .i(_91[3:1]), .done_(_91[0:0]) );
    assign _1660 = _91[0:0];

    /* aliases */
    assign data_0 = data;
    assign data_2 = data_1;
    assign data_4 = data_3;
    assign data_5 = data_3;
    assign data_6 = data_3;
    assign data_8 = data_7;
    assign data_9 = data_7;
    assign data_10 = data_7;
    assign data_12 = data_11;
    assign data_14 = data_13;
    assign data_16 = data_15;
    assign data_17 = data_15;
    assign data_18 = data_15;
    assign data_20 = data_19;
    assign data_21 = data_19;
    assign data_22 = data_19;
    assign data_24 = data_23;
    assign data_26 = data_25;
    assign data_28 = data_27;
    assign data_29 = data_27;
    assign data_30 = data_27;
    assign data_32 = data_31;
    assign data_33 = data_31;
    assign data_34 = data_31;
    assign data_36 = data_35;
    assign data_38 = data_37;
    assign data_40 = data_39;
    assign data_41 = data_39;
    assign data_42 = data_39;
    assign data_44 = data_43;
    assign data_45 = data_43;
    assign data_46 = data_43;
    assign data_48 = data_47;
    assign data_50 = data_49;
    assign data_52 = data_51;
    assign data_53 = data_51;
    assign data_54 = data_51;
    assign data_56 = data_55;
    assign data_57 = data_55;
    assign data_58 = data_55;
    assign data_60 = data_59;
    assign data_62 = data_61;
    assign data_64 = data_63;
    assign data_65 = data_63;
    assign data_66 = data_63;
    assign data_68 = data_67;
    assign data_69 = data_67;
    assign data_70 = data_67;
    assign data_72 = data_71;
    assign data_74 = data_73;
    assign data_76 = data_75;
    assign data_77 = data_75;
    assign data_78 = data_75;
    assign data_80 = data_79;
    assign data_81 = data_79;
    assign data_82 = data_79;
    assign data_84 = data_83;
    assign data_86 = data_85;
    assign data_88 = data_87;
    assign data_89 = data_87;
    assign data_90 = data_87;
    assign data_92 = data_91;
    assign data_93 = data_91;
    assign data_94 = data_91;

    /* output assignments */
    assign done_ = _1660;
    assign rd_q0 = _1659;
    assign rd_q1 = _1475;
    assign rd_q2 = _1291;
    assign rd_q3 = _1107;
    assign rd_q4 = _923;
    assign rd_q5 = _739;
    assign rd_q6 = _555;
    assign rd_q7 = _371;

endmodule
module dp_23 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0010110101010100000011011110111011010110010100110001101011101000;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0010101001011001010100000010000110010000100101110100011001111101;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0101101010011100111100001000011100111110010010010000110000101110;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1010001101110111101111000010110101111101000101111110101011000110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0000001111101000110111111101001001001110100011100111100000011111;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1011101000100101111010110101110011010001100101110000101011101011;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_24 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0011111001001010001001101011111101110010010000001011101010111010;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0011000010100101000101000101111001000110100000100110000111011001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0110011101011010100011100010100100001000011111001101101001001010;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0000101111111101100110101110100101111000100111010010010010100100;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0000001001111011000100111011001010010011010011011101111001111100;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1111111101011100001000000110011010110000001001110010101101001011;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0100000000001010011100001110010111000101111110001100111000110011;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_25 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0111010100110110111000101101011010010001100100010001111101010110;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0000110011000010001010101100101000000111101110001000000000100010;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0111001000110011101111100110101010100000101011000011100010011000;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0101001001010011010110011100100111011110000001110100111001010010;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1010000011011100010101000100001100110010011011110100111011000101;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0101110010000010010001101000010101000000100001101011001000100011;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0000011100001011110100010000110110100011110110100100101101101110;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_26 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1110101110110100001110011000001101010010101110001110101101001001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0100001101001001101100101111100001110111000100100000100100101110;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0111001001000001100001111101100111010000000111101110111101101001;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1010100110001010110101010011000100100110101001101111101110101001;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0110101111001100100110001011001000101110101111101111010110101001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0111010010100011111001001101111110000010101010011101010011011100;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0101001110100110001000001111011110000111100111011011010111100001;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_27 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1010010011111010110011100011111011010001110100111011000111100110;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0010110101010100000011011110111011010110010100110001101011101000;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0100101111010011001001111101111001111010100010111010100101011100;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0011101110101011111110001010011100001011100100000001011011010111;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0011001010101001010101000011100000101111110100000000100010101001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1001010110000011011011011110011100001111001100011100101111111010;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0101010011010111101011100001010011111111011110000011001100001001;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_28 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0111011110011110111111110110000011000011011101000101101100101101;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1000100001000000000010001010111011110000011011011110010100110100;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0100010111000111001011011001011100011001101100111010011010110011;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1000010001111100010101000001111110111110110111001011110100110010;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0110010011100110000100100001110100111010001101101101000100011110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1100000100011100001110111010011001111110100101100110010100000101;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0100110100101011001101101011101110010010101100011011100111111010;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_29 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0111111011110111100011010110100101100101011001110101010011100001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1010110010001000101010001101111011000001110101011110111111011111;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0011000010100101000101000101111001000110100000100110000111011001;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0101101010011100111100001000011100111110010010010000110000101110;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0111001100001110001111011101000101111010000101110111100100101011;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0011100110101111101011010110110000110010100010110001011011110110;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0000001101001101110010111010010110001010110001010000000000111110;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_30 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _231 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _230 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _229 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _228 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _227 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _226 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1110001100111111001111111001011100111001101010000000000101001111;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1001100101000001000011111011100001010111110101010010000001011011;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0110110101111000001010110001011000001010010010011101111000011001;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0001110101100010001100010001100100101000001010010100100111001010;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1110111001111000010110101100100001101010011001001010001000010001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1010011001111001100010101011001010101101111110001111101110010010;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0111000100111110100110011110111110011000000010111100110110100000;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module parallel_cores_2 (
    wr_d7,
    wr_d6,
    wr_d5,
    wr_d4,
    wr_d3,
    wr_d2,
    wr_d1,
    wr_d0,
    wr_addr,
    wr_en,
    rd_addr,
    rd_en,
    flip,
    first_4step_pass,
    first_iter,
    start,
    clear,
    clock,
    done_,
    rd_q0,
    rd_q1,
    rd_q2,
    rd_q3,
    rd_q4,
    rd_q5,
    rd_q6,
    rd_q7
);

    input [63:0] wr_d7;
    input [63:0] wr_d6;
    input [63:0] wr_d5;
    input [63:0] wr_d4;
    input [63:0] wr_d3;
    input [63:0] wr_d2;
    input [63:0] wr_d1;
    input [63:0] wr_d0;
    input [5:0] wr_addr;
    input [7:0] wr_en;
    input [5:0] rd_addr;
    input [7:0] rd_en;
    input flip;
    input first_4step_pass;
    input first_iter;
    input start;
    input clear;
    input clock;
    output done_;
    output [63:0] rd_q0;
    output [63:0] rd_q1;
    output [63:0] rd_q2;
    output [63:0] rd_q3;
    output [63:0] rd_q4;
    output [63:0] rd_q5;
    output [63:0] rd_q6;
    output [63:0] rd_q7;

    /* signal declarations */
    wire [5:0] address;
    wire write_enable;
    wire [5:0] address_0;
    wire _362;
    wire read_enable;
    wire _360;
    wire write_enable_0;
    wire _364;
    wire [131:0] _369;
    wire [63:0] _370;
    wire [5:0] _355 = 6'b000000;
    wire [5:0] address_1;
    wire _353;
    wire write_enable_1;
    wire [63:0] _267;
    wire [63:0] _266;
    wire [63:0] _268;
    wire [63:0] _264;
    wire [63:0] _263;
    wire [63:0] q1;
    wire [63:0] _269;
    wire [5:0] address_2;
    wire write_enable_2 = 1'b0;
    wire _254;
    wire read_enable_0;
    wire [5:0] address_3;
    wire _250;
    wire read_enable_1;
    wire _248;
    wire write_enable_3;
    wire _252;
    wire [131:0] _259;
    wire [63:0] _260;
    wire [63:0] data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_0;
    wire [5:0] _242 = 6'b000000;
    wire _240;
    wire _239;
    wire _238;
    wire _237;
    wire _236;
    wire _235;
    wire [5:0] _241;
    wire [5:0] address_4;
    wire write_enable_4 = 1'b0;
    wire _232;
    wire read_enable_2;
    wire [63:0] data_1;
    wire [63:0] data_2;
    wire _229;
    wire _228;
    wire _227;
    wire _226;
    wire _225;
    wire _224;
    wire [5:0] _230;
    wire [5:0] address_5;
    wire _221;
    wire read_enable_3;
    wire _219;
    wire write_enable_5;
    wire _223;
    wire [131:0] _246;
    wire [63:0] _247;
    wire _87 = 1'b0;
    wire _86 = 1'b0;
    wire _89;
    wire _3;
    reg PHASE;
    wire [63:0] _261;
    wire [5:0] address_6;
    wire _211;
    wire read_enable_4;
    wire write_enable_6;
    wire _213;
    wire [5:0] address_7;
    wire _206;
    wire read_enable_5;
    wire _204;
    wire write_enable_7;
    wire _208;
    wire [131:0] _216;
    wire [63:0] _217;
    wire [63:0] _283;
    wire [63:0] data_3;
    wire [63:0] data_4;
    wire [63:0] data_5;
    wire [63:0] data_6;
    wire [5:0] address_8;
    wire _169;
    wire read_enable_6;
    wire _166;
    wire _167;
    wire write_enable_8;
    wire _171;
    wire [5:0] address_9;
    wire _134;
    wire read_enable_7;
    wire _131;
    wire _132;
    wire write_enable_9;
    wire _136;
    wire [131:0] _202;
    wire [63:0] _203;
    wire _98 = 1'b0;
    wire _97 = 1'b0;
    wire _284;
    wire _5;
    reg PHASE_0;
    wire [63:0] q0;
    wire _94 = 1'b0;
    wire _93 = 1'b0;
    reg _96;
    wire [63:0] _262;
    wire [191:0] _282;
    wire [63:0] _285;
    wire [63:0] data_7;
    wire [63:0] data_8;
    wire [63:0] data_9;
    wire [63:0] data_10;
    wire [5:0] address_10;
    wire _349;
    wire _348;
    wire read_enable_8;
    wire _342 = 1'b0;
    wire _341 = 1'b0;
    wire _339 = 1'b0;
    wire _338 = 1'b0;
    wire _336 = 1'b0;
    wire _335 = 1'b0;
    wire _333 = 1'b0;
    wire _332 = 1'b0;
    wire _330 = 1'b0;
    wire _329 = 1'b0;
    wire _327 = 1'b0;
    wire _326 = 1'b0;
    wire _324 = 1'b0;
    wire _323 = 1'b0;
    wire _321 = 1'b0;
    wire _320 = 1'b0;
    wire _318 = 1'b0;
    wire _317 = 1'b0;
    reg _319;
    reg _322;
    reg _325;
    reg _328;
    reg _331;
    reg _334;
    reg _337;
    reg _340;
    reg _343;
    wire _344;
    wire _315 = 1'b0;
    wire _314 = 1'b0;
    wire _312 = 1'b0;
    wire _311 = 1'b0;
    wire _309 = 1'b0;
    wire _308 = 1'b0;
    wire _306 = 1'b0;
    wire _305 = 1'b0;
    wire _303 = 1'b0;
    wire _302 = 1'b0;
    wire _300 = 1'b0;
    wire _299 = 1'b0;
    wire _297 = 1'b0;
    wire _296 = 1'b0;
    wire _294 = 1'b0;
    wire _293 = 1'b0;
    wire _291 = 1'b0;
    wire _290 = 1'b0;
    reg _292;
    reg _295;
    reg _298;
    reg _301;
    reg _304;
    reg _307;
    reg _310;
    reg _313;
    reg _316;
    wire _345;
    wire _346;
    wire write_enable_10;
    wire _351;
    wire [131:0] _358;
    wire [63:0] _359;
    wire _287 = 1'b0;
    wire _286 = 1'b0;
    wire _289;
    wire _7;
    reg PHASE_1;
    wire [63:0] _371;
    wire [5:0] address_11;
    wire write_enable_11;
    wire [5:0] address_12;
    wire _546;
    wire read_enable_9;
    wire _544;
    wire write_enable_12;
    wire _548;
    wire [131:0] _553;
    wire [63:0] _554;
    wire [5:0] _539 = 6'b000000;
    wire [5:0] address_13;
    wire _537;
    wire write_enable_13;
    wire [63:0] _462;
    wire [63:0] _461;
    wire [63:0] _463;
    wire [63:0] _459;
    wire [63:0] _458;
    wire [63:0] q1_0;
    wire [63:0] _464;
    wire [5:0] address_14;
    wire write_enable_14 = 1'b0;
    wire _449;
    wire read_enable_10;
    wire [5:0] address_15;
    wire _445;
    wire read_enable_11;
    wire _443;
    wire write_enable_15;
    wire _447;
    wire [131:0] _454;
    wire [63:0] _455;
    wire [63:0] data_11 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_12;
    wire [5:0] _437 = 6'b000000;
    wire _435;
    wire _434;
    wire _433;
    wire _432;
    wire _431;
    wire _430;
    wire [5:0] _436;
    wire [5:0] address_16;
    wire write_enable_16 = 1'b0;
    wire _427;
    wire read_enable_12;
    wire [63:0] data_13;
    wire [63:0] data_14;
    wire _424;
    wire _423;
    wire _422;
    wire _421;
    wire _420;
    wire _419;
    wire [5:0] _425;
    wire [5:0] address_17;
    wire _416;
    wire read_enable_13;
    wire _414;
    wire write_enable_17;
    wire _418;
    wire [131:0] _441;
    wire [63:0] _442;
    wire _373 = 1'b0;
    wire _372 = 1'b0;
    wire _375;
    wire _11;
    reg PHASE_2;
    wire [63:0] _456;
    wire [5:0] address_18;
    wire _406;
    wire read_enable_14;
    wire write_enable_18;
    wire _408;
    wire [5:0] address_19;
    wire _401;
    wire read_enable_15;
    wire _399;
    wire write_enable_19;
    wire _403;
    wire [131:0] _411;
    wire [63:0] _412;
    wire [63:0] _467;
    wire [63:0] data_15;
    wire [63:0] data_16;
    wire [63:0] data_17;
    wire [63:0] data_18;
    wire [5:0] address_20;
    wire _392;
    wire read_enable_16;
    wire _389;
    wire _390;
    wire write_enable_20;
    wire _394;
    wire [5:0] address_21;
    wire _385;
    wire read_enable_17;
    wire _382;
    wire _383;
    wire write_enable_21;
    wire _387;
    wire [131:0] _397;
    wire [63:0] _398;
    wire _380 = 1'b0;
    wire _379 = 1'b0;
    wire _468;
    wire _13;
    reg PHASE_3;
    wire [63:0] q0_0;
    wire _377 = 1'b0;
    wire _376 = 1'b0;
    reg _378;
    wire [63:0] _457;
    wire [191:0] _466;
    wire [63:0] _469;
    wire [63:0] data_19;
    wire [63:0] data_20;
    wire [63:0] data_21;
    wire [63:0] data_22;
    wire [5:0] address_22;
    wire _533;
    wire _532;
    wire read_enable_18;
    wire _526 = 1'b0;
    wire _525 = 1'b0;
    wire _523 = 1'b0;
    wire _522 = 1'b0;
    wire _520 = 1'b0;
    wire _519 = 1'b0;
    wire _517 = 1'b0;
    wire _516 = 1'b0;
    wire _514 = 1'b0;
    wire _513 = 1'b0;
    wire _511 = 1'b0;
    wire _510 = 1'b0;
    wire _508 = 1'b0;
    wire _507 = 1'b0;
    wire _505 = 1'b0;
    wire _504 = 1'b0;
    wire _502 = 1'b0;
    wire _501 = 1'b0;
    reg _503;
    reg _506;
    reg _509;
    reg _512;
    reg _515;
    reg _518;
    reg _521;
    reg _524;
    reg _527;
    wire _528;
    wire _499 = 1'b0;
    wire _498 = 1'b0;
    wire _496 = 1'b0;
    wire _495 = 1'b0;
    wire _493 = 1'b0;
    wire _492 = 1'b0;
    wire _490 = 1'b0;
    wire _489 = 1'b0;
    wire _487 = 1'b0;
    wire _486 = 1'b0;
    wire _484 = 1'b0;
    wire _483 = 1'b0;
    wire _481 = 1'b0;
    wire _480 = 1'b0;
    wire _478 = 1'b0;
    wire _477 = 1'b0;
    wire _475 = 1'b0;
    wire _474 = 1'b0;
    reg _476;
    reg _479;
    reg _482;
    reg _485;
    reg _488;
    reg _491;
    reg _494;
    reg _497;
    reg _500;
    wire _529;
    wire _530;
    wire write_enable_22;
    wire _535;
    wire [131:0] _542;
    wire [63:0] _543;
    wire _471 = 1'b0;
    wire _470 = 1'b0;
    wire _473;
    wire _15;
    reg PHASE_4;
    wire [63:0] _555;
    wire [5:0] address_23;
    wire write_enable_23;
    wire [5:0] address_24;
    wire _730;
    wire read_enable_19;
    wire _728;
    wire write_enable_24;
    wire _732;
    wire [131:0] _737;
    wire [63:0] _738;
    wire [5:0] _723 = 6'b000000;
    wire [5:0] address_25;
    wire _721;
    wire write_enable_25;
    wire [63:0] _646;
    wire [63:0] _645;
    wire [63:0] _647;
    wire [63:0] _643;
    wire [63:0] _642;
    wire [63:0] q1_1;
    wire [63:0] _648;
    wire [5:0] address_26;
    wire write_enable_26 = 1'b0;
    wire _633;
    wire read_enable_20;
    wire [5:0] address_27;
    wire _629;
    wire read_enable_21;
    wire _627;
    wire write_enable_27;
    wire _631;
    wire [131:0] _638;
    wire [63:0] _639;
    wire [63:0] data_23 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_24;
    wire [5:0] _621 = 6'b000000;
    wire _619;
    wire _618;
    wire _617;
    wire _616;
    wire _615;
    wire _614;
    wire [5:0] _620;
    wire [5:0] address_28;
    wire write_enable_28 = 1'b0;
    wire _611;
    wire read_enable_22;
    wire [63:0] data_25;
    wire [63:0] data_26;
    wire _608;
    wire _607;
    wire _606;
    wire _605;
    wire _604;
    wire _603;
    wire [5:0] _609;
    wire [5:0] address_29;
    wire _600;
    wire read_enable_23;
    wire _598;
    wire write_enable_29;
    wire _602;
    wire [131:0] _625;
    wire [63:0] _626;
    wire _557 = 1'b0;
    wire _556 = 1'b0;
    wire _559;
    wire _19;
    reg PHASE_5;
    wire [63:0] _640;
    wire [5:0] address_30;
    wire _590;
    wire read_enable_24;
    wire write_enable_30;
    wire _592;
    wire [5:0] address_31;
    wire _585;
    wire read_enable_25;
    wire _583;
    wire write_enable_31;
    wire _587;
    wire [131:0] _595;
    wire [63:0] _596;
    wire [63:0] _651;
    wire [63:0] data_27;
    wire [63:0] data_28;
    wire [63:0] data_29;
    wire [63:0] data_30;
    wire [5:0] address_32;
    wire _576;
    wire read_enable_26;
    wire _573;
    wire _574;
    wire write_enable_32;
    wire _578;
    wire [5:0] address_33;
    wire _569;
    wire read_enable_27;
    wire _566;
    wire _567;
    wire write_enable_33;
    wire _571;
    wire [131:0] _581;
    wire [63:0] _582;
    wire _564 = 1'b0;
    wire _563 = 1'b0;
    wire _652;
    wire _21;
    reg PHASE_6;
    wire [63:0] q0_1;
    wire _561 = 1'b0;
    wire _560 = 1'b0;
    reg _562;
    wire [63:0] _641;
    wire [191:0] _650;
    wire [63:0] _653;
    wire [63:0] data_31;
    wire [63:0] data_32;
    wire [63:0] data_33;
    wire [63:0] data_34;
    wire [5:0] address_34;
    wire _717;
    wire _716;
    wire read_enable_28;
    wire _710 = 1'b0;
    wire _709 = 1'b0;
    wire _707 = 1'b0;
    wire _706 = 1'b0;
    wire _704 = 1'b0;
    wire _703 = 1'b0;
    wire _701 = 1'b0;
    wire _700 = 1'b0;
    wire _698 = 1'b0;
    wire _697 = 1'b0;
    wire _695 = 1'b0;
    wire _694 = 1'b0;
    wire _692 = 1'b0;
    wire _691 = 1'b0;
    wire _689 = 1'b0;
    wire _688 = 1'b0;
    wire _686 = 1'b0;
    wire _685 = 1'b0;
    reg _687;
    reg _690;
    reg _693;
    reg _696;
    reg _699;
    reg _702;
    reg _705;
    reg _708;
    reg _711;
    wire _712;
    wire _683 = 1'b0;
    wire _682 = 1'b0;
    wire _680 = 1'b0;
    wire _679 = 1'b0;
    wire _677 = 1'b0;
    wire _676 = 1'b0;
    wire _674 = 1'b0;
    wire _673 = 1'b0;
    wire _671 = 1'b0;
    wire _670 = 1'b0;
    wire _668 = 1'b0;
    wire _667 = 1'b0;
    wire _665 = 1'b0;
    wire _664 = 1'b0;
    wire _662 = 1'b0;
    wire _661 = 1'b0;
    wire _659 = 1'b0;
    wire _658 = 1'b0;
    reg _660;
    reg _663;
    reg _666;
    reg _669;
    reg _672;
    reg _675;
    reg _678;
    reg _681;
    reg _684;
    wire _713;
    wire _714;
    wire write_enable_34;
    wire _719;
    wire [131:0] _726;
    wire [63:0] _727;
    wire _655 = 1'b0;
    wire _654 = 1'b0;
    wire _657;
    wire _23;
    reg PHASE_7;
    wire [63:0] _739;
    wire [5:0] address_35;
    wire write_enable_35;
    wire [5:0] address_36;
    wire _914;
    wire read_enable_29;
    wire _912;
    wire write_enable_36;
    wire _916;
    wire [131:0] _921;
    wire [63:0] _922;
    wire [5:0] _907 = 6'b000000;
    wire [5:0] address_37;
    wire _905;
    wire write_enable_37;
    wire [63:0] _830;
    wire [63:0] _829;
    wire [63:0] _831;
    wire [63:0] _827;
    wire [63:0] _826;
    wire [63:0] q1_2;
    wire [63:0] _832;
    wire [5:0] address_38;
    wire write_enable_38 = 1'b0;
    wire _817;
    wire read_enable_30;
    wire [5:0] address_39;
    wire _813;
    wire read_enable_31;
    wire _811;
    wire write_enable_39;
    wire _815;
    wire [131:0] _822;
    wire [63:0] _823;
    wire [63:0] data_35 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_36;
    wire [5:0] _805 = 6'b000000;
    wire _803;
    wire _802;
    wire _801;
    wire _800;
    wire _799;
    wire _798;
    wire [5:0] _804;
    wire [5:0] address_40;
    wire write_enable_40 = 1'b0;
    wire _795;
    wire read_enable_32;
    wire [63:0] data_37;
    wire [63:0] data_38;
    wire _792;
    wire _791;
    wire _790;
    wire _789;
    wire _788;
    wire _787;
    wire [5:0] _793;
    wire [5:0] address_41;
    wire _784;
    wire read_enable_33;
    wire _782;
    wire write_enable_41;
    wire _786;
    wire [131:0] _809;
    wire [63:0] _810;
    wire _741 = 1'b0;
    wire _740 = 1'b0;
    wire _743;
    wire _27;
    reg PHASE_8;
    wire [63:0] _824;
    wire [5:0] address_42;
    wire _774;
    wire read_enable_34;
    wire write_enable_42;
    wire _776;
    wire [5:0] address_43;
    wire _769;
    wire read_enable_35;
    wire _767;
    wire write_enable_43;
    wire _771;
    wire [131:0] _779;
    wire [63:0] _780;
    wire [63:0] _835;
    wire [63:0] data_39;
    wire [63:0] data_40;
    wire [63:0] data_41;
    wire [63:0] data_42;
    wire [5:0] address_44;
    wire _760;
    wire read_enable_36;
    wire _757;
    wire _758;
    wire write_enable_44;
    wire _762;
    wire [5:0] address_45;
    wire _753;
    wire read_enable_37;
    wire _750;
    wire _751;
    wire write_enable_45;
    wire _755;
    wire [131:0] _765;
    wire [63:0] _766;
    wire _748 = 1'b0;
    wire _747 = 1'b0;
    wire _836;
    wire _29;
    reg PHASE_9;
    wire [63:0] q0_2;
    wire _745 = 1'b0;
    wire _744 = 1'b0;
    reg _746;
    wire [63:0] _825;
    wire [191:0] _834;
    wire [63:0] _837;
    wire [63:0] data_43;
    wire [63:0] data_44;
    wire [63:0] data_45;
    wire [63:0] data_46;
    wire [5:0] address_46;
    wire _901;
    wire _900;
    wire read_enable_38;
    wire _894 = 1'b0;
    wire _893 = 1'b0;
    wire _891 = 1'b0;
    wire _890 = 1'b0;
    wire _888 = 1'b0;
    wire _887 = 1'b0;
    wire _885 = 1'b0;
    wire _884 = 1'b0;
    wire _882 = 1'b0;
    wire _881 = 1'b0;
    wire _879 = 1'b0;
    wire _878 = 1'b0;
    wire _876 = 1'b0;
    wire _875 = 1'b0;
    wire _873 = 1'b0;
    wire _872 = 1'b0;
    wire _870 = 1'b0;
    wire _869 = 1'b0;
    reg _871;
    reg _874;
    reg _877;
    reg _880;
    reg _883;
    reg _886;
    reg _889;
    reg _892;
    reg _895;
    wire _896;
    wire _867 = 1'b0;
    wire _866 = 1'b0;
    wire _864 = 1'b0;
    wire _863 = 1'b0;
    wire _861 = 1'b0;
    wire _860 = 1'b0;
    wire _858 = 1'b0;
    wire _857 = 1'b0;
    wire _855 = 1'b0;
    wire _854 = 1'b0;
    wire _852 = 1'b0;
    wire _851 = 1'b0;
    wire _849 = 1'b0;
    wire _848 = 1'b0;
    wire _846 = 1'b0;
    wire _845 = 1'b0;
    wire _843 = 1'b0;
    wire _842 = 1'b0;
    reg _844;
    reg _847;
    reg _850;
    reg _853;
    reg _856;
    reg _859;
    reg _862;
    reg _865;
    reg _868;
    wire _897;
    wire _898;
    wire write_enable_46;
    wire _903;
    wire [131:0] _910;
    wire [63:0] _911;
    wire _839 = 1'b0;
    wire _838 = 1'b0;
    wire _841;
    wire _31;
    reg PHASE_10;
    wire [63:0] _923;
    wire [5:0] address_47;
    wire write_enable_47;
    wire [5:0] address_48;
    wire _1098;
    wire read_enable_39;
    wire _1096;
    wire write_enable_48;
    wire _1100;
    wire [131:0] _1105;
    wire [63:0] _1106;
    wire [5:0] _1091 = 6'b000000;
    wire [5:0] address_49;
    wire _1089;
    wire write_enable_49;
    wire [63:0] _1014;
    wire [63:0] _1013;
    wire [63:0] _1015;
    wire [63:0] _1011;
    wire [63:0] _1010;
    wire [63:0] q1_3;
    wire [63:0] _1016;
    wire [5:0] address_50;
    wire write_enable_50 = 1'b0;
    wire _1001;
    wire read_enable_40;
    wire [5:0] address_51;
    wire _997;
    wire read_enable_41;
    wire _995;
    wire write_enable_51;
    wire _999;
    wire [131:0] _1006;
    wire [63:0] _1007;
    wire [63:0] data_47 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_48;
    wire [5:0] _989 = 6'b000000;
    wire _987;
    wire _986;
    wire _985;
    wire _984;
    wire _983;
    wire _982;
    wire [5:0] _988;
    wire [5:0] address_52;
    wire write_enable_52 = 1'b0;
    wire _979;
    wire read_enable_42;
    wire [63:0] data_49;
    wire [63:0] data_50;
    wire _976;
    wire _975;
    wire _974;
    wire _973;
    wire _972;
    wire _971;
    wire [5:0] _977;
    wire [5:0] address_53;
    wire _968;
    wire read_enable_43;
    wire _966;
    wire write_enable_53;
    wire _970;
    wire [131:0] _993;
    wire [63:0] _994;
    wire _925 = 1'b0;
    wire _924 = 1'b0;
    wire _927;
    wire _35;
    reg PHASE_11;
    wire [63:0] _1008;
    wire [5:0] address_54;
    wire _958;
    wire read_enable_44;
    wire write_enable_54;
    wire _960;
    wire [5:0] address_55;
    wire _953;
    wire read_enable_45;
    wire _951;
    wire write_enable_55;
    wire _955;
    wire [131:0] _963;
    wire [63:0] _964;
    wire [63:0] _1019;
    wire [63:0] data_51;
    wire [63:0] data_52;
    wire [63:0] data_53;
    wire [63:0] data_54;
    wire [5:0] address_56;
    wire _944;
    wire read_enable_46;
    wire _941;
    wire _942;
    wire write_enable_56;
    wire _946;
    wire [5:0] address_57;
    wire _937;
    wire read_enable_47;
    wire _934;
    wire _935;
    wire write_enable_57;
    wire _939;
    wire [131:0] _949;
    wire [63:0] _950;
    wire _932 = 1'b0;
    wire _931 = 1'b0;
    wire _1020;
    wire _37;
    reg PHASE_12;
    wire [63:0] q0_3;
    wire _929 = 1'b0;
    wire _928 = 1'b0;
    reg _930;
    wire [63:0] _1009;
    wire [191:0] _1018;
    wire [63:0] _1021;
    wire [63:0] data_55;
    wire [63:0] data_56;
    wire [63:0] data_57;
    wire [63:0] data_58;
    wire [5:0] address_58;
    wire _1085;
    wire _1084;
    wire read_enable_48;
    wire _1078 = 1'b0;
    wire _1077 = 1'b0;
    wire _1075 = 1'b0;
    wire _1074 = 1'b0;
    wire _1072 = 1'b0;
    wire _1071 = 1'b0;
    wire _1069 = 1'b0;
    wire _1068 = 1'b0;
    wire _1066 = 1'b0;
    wire _1065 = 1'b0;
    wire _1063 = 1'b0;
    wire _1062 = 1'b0;
    wire _1060 = 1'b0;
    wire _1059 = 1'b0;
    wire _1057 = 1'b0;
    wire _1056 = 1'b0;
    wire _1054 = 1'b0;
    wire _1053 = 1'b0;
    reg _1055;
    reg _1058;
    reg _1061;
    reg _1064;
    reg _1067;
    reg _1070;
    reg _1073;
    reg _1076;
    reg _1079;
    wire _1080;
    wire _1051 = 1'b0;
    wire _1050 = 1'b0;
    wire _1048 = 1'b0;
    wire _1047 = 1'b0;
    wire _1045 = 1'b0;
    wire _1044 = 1'b0;
    wire _1042 = 1'b0;
    wire _1041 = 1'b0;
    wire _1039 = 1'b0;
    wire _1038 = 1'b0;
    wire _1036 = 1'b0;
    wire _1035 = 1'b0;
    wire _1033 = 1'b0;
    wire _1032 = 1'b0;
    wire _1030 = 1'b0;
    wire _1029 = 1'b0;
    wire _1027 = 1'b0;
    wire _1026 = 1'b0;
    reg _1028;
    reg _1031;
    reg _1034;
    reg _1037;
    reg _1040;
    reg _1043;
    reg _1046;
    reg _1049;
    reg _1052;
    wire _1081;
    wire _1082;
    wire write_enable_58;
    wire _1087;
    wire [131:0] _1094;
    wire [63:0] _1095;
    wire _1023 = 1'b0;
    wire _1022 = 1'b0;
    wire _1025;
    wire _39;
    reg PHASE_13;
    wire [63:0] _1107;
    wire [5:0] address_59;
    wire write_enable_59;
    wire [5:0] address_60;
    wire _1282;
    wire read_enable_49;
    wire _1280;
    wire write_enable_60;
    wire _1284;
    wire [131:0] _1289;
    wire [63:0] _1290;
    wire [5:0] _1275 = 6'b000000;
    wire [5:0] address_61;
    wire _1273;
    wire write_enable_61;
    wire [63:0] _1198;
    wire [63:0] _1197;
    wire [63:0] _1199;
    wire [63:0] _1195;
    wire [63:0] _1194;
    wire [63:0] q1_4;
    wire [63:0] _1200;
    wire [5:0] address_62;
    wire write_enable_62 = 1'b0;
    wire _1185;
    wire read_enable_50;
    wire [5:0] address_63;
    wire _1181;
    wire read_enable_51;
    wire _1179;
    wire write_enable_63;
    wire _1183;
    wire [131:0] _1190;
    wire [63:0] _1191;
    wire [63:0] data_59 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_60;
    wire [5:0] _1173 = 6'b000000;
    wire _1171;
    wire _1170;
    wire _1169;
    wire _1168;
    wire _1167;
    wire _1166;
    wire [5:0] _1172;
    wire [5:0] address_64;
    wire write_enable_64 = 1'b0;
    wire _1163;
    wire read_enable_52;
    wire [63:0] data_61;
    wire [63:0] data_62;
    wire _1160;
    wire _1159;
    wire _1158;
    wire _1157;
    wire _1156;
    wire _1155;
    wire [5:0] _1161;
    wire [5:0] address_65;
    wire _1152;
    wire read_enable_53;
    wire _1150;
    wire write_enable_65;
    wire _1154;
    wire [131:0] _1177;
    wire [63:0] _1178;
    wire _1109 = 1'b0;
    wire _1108 = 1'b0;
    wire _1111;
    wire _43;
    reg PHASE_14;
    wire [63:0] _1192;
    wire [5:0] address_66;
    wire _1142;
    wire read_enable_54;
    wire write_enable_66;
    wire _1144;
    wire [5:0] address_67;
    wire _1137;
    wire read_enable_55;
    wire _1135;
    wire write_enable_67;
    wire _1139;
    wire [131:0] _1147;
    wire [63:0] _1148;
    wire [63:0] _1203;
    wire [63:0] data_63;
    wire [63:0] data_64;
    wire [63:0] data_65;
    wire [63:0] data_66;
    wire [5:0] address_68;
    wire _1128;
    wire read_enable_56;
    wire _1125;
    wire _1126;
    wire write_enable_68;
    wire _1130;
    wire [5:0] address_69;
    wire _1121;
    wire read_enable_57;
    wire _1118;
    wire _1119;
    wire write_enable_69;
    wire _1123;
    wire [131:0] _1133;
    wire [63:0] _1134;
    wire _1116 = 1'b0;
    wire _1115 = 1'b0;
    wire _1204;
    wire _45;
    reg PHASE_15;
    wire [63:0] q0_4;
    wire _1113 = 1'b0;
    wire _1112 = 1'b0;
    reg _1114;
    wire [63:0] _1193;
    wire [191:0] _1202;
    wire [63:0] _1205;
    wire [63:0] data_67;
    wire [63:0] data_68;
    wire [63:0] data_69;
    wire [63:0] data_70;
    wire [5:0] address_70;
    wire _1269;
    wire _1268;
    wire read_enable_58;
    wire _1262 = 1'b0;
    wire _1261 = 1'b0;
    wire _1259 = 1'b0;
    wire _1258 = 1'b0;
    wire _1256 = 1'b0;
    wire _1255 = 1'b0;
    wire _1253 = 1'b0;
    wire _1252 = 1'b0;
    wire _1250 = 1'b0;
    wire _1249 = 1'b0;
    wire _1247 = 1'b0;
    wire _1246 = 1'b0;
    wire _1244 = 1'b0;
    wire _1243 = 1'b0;
    wire _1241 = 1'b0;
    wire _1240 = 1'b0;
    wire _1238 = 1'b0;
    wire _1237 = 1'b0;
    reg _1239;
    reg _1242;
    reg _1245;
    reg _1248;
    reg _1251;
    reg _1254;
    reg _1257;
    reg _1260;
    reg _1263;
    wire _1264;
    wire _1235 = 1'b0;
    wire _1234 = 1'b0;
    wire _1232 = 1'b0;
    wire _1231 = 1'b0;
    wire _1229 = 1'b0;
    wire _1228 = 1'b0;
    wire _1226 = 1'b0;
    wire _1225 = 1'b0;
    wire _1223 = 1'b0;
    wire _1222 = 1'b0;
    wire _1220 = 1'b0;
    wire _1219 = 1'b0;
    wire _1217 = 1'b0;
    wire _1216 = 1'b0;
    wire _1214 = 1'b0;
    wire _1213 = 1'b0;
    wire _1211 = 1'b0;
    wire _1210 = 1'b0;
    reg _1212;
    reg _1215;
    reg _1218;
    reg _1221;
    reg _1224;
    reg _1227;
    reg _1230;
    reg _1233;
    reg _1236;
    wire _1265;
    wire _1266;
    wire write_enable_70;
    wire _1271;
    wire [131:0] _1278;
    wire [63:0] _1279;
    wire _1207 = 1'b0;
    wire _1206 = 1'b0;
    wire _1209;
    wire _47;
    reg PHASE_16;
    wire [63:0] _1291;
    wire [5:0] address_71;
    wire write_enable_71;
    wire [5:0] address_72;
    wire _1466;
    wire read_enable_59;
    wire _1464;
    wire write_enable_72;
    wire _1468;
    wire [131:0] _1473;
    wire [63:0] _1474;
    wire [5:0] _1459 = 6'b000000;
    wire [5:0] address_73;
    wire _1457;
    wire write_enable_73;
    wire [63:0] _1382;
    wire [63:0] _1381;
    wire [63:0] _1383;
    wire [63:0] _1379;
    wire [63:0] _1378;
    wire [63:0] q1_5;
    wire [63:0] _1384;
    wire [5:0] address_74;
    wire write_enable_74 = 1'b0;
    wire _1369;
    wire read_enable_60;
    wire [5:0] address_75;
    wire _1365;
    wire read_enable_61;
    wire _1363;
    wire write_enable_75;
    wire _1367;
    wire [131:0] _1374;
    wire [63:0] _1375;
    wire [63:0] data_71 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_72;
    wire [5:0] _1357 = 6'b000000;
    wire _1355;
    wire _1354;
    wire _1353;
    wire _1352;
    wire _1351;
    wire _1350;
    wire [5:0] _1356;
    wire [5:0] address_76;
    wire write_enable_76 = 1'b0;
    wire _1347;
    wire read_enable_62;
    wire [63:0] data_73;
    wire [63:0] data_74;
    wire _1344;
    wire _1343;
    wire _1342;
    wire _1341;
    wire _1340;
    wire _1339;
    wire [5:0] _1345;
    wire [5:0] address_77;
    wire _1336;
    wire read_enable_63;
    wire _1334;
    wire write_enable_77;
    wire _1338;
    wire [131:0] _1361;
    wire [63:0] _1362;
    wire _1293 = 1'b0;
    wire _1292 = 1'b0;
    wire _1295;
    wire _51;
    reg PHASE_17;
    wire [63:0] _1376;
    wire [5:0] address_78;
    wire _1326;
    wire read_enable_64;
    wire write_enable_78;
    wire _1328;
    wire [5:0] address_79;
    wire _1321;
    wire read_enable_65;
    wire _1319;
    wire write_enable_79;
    wire _1323;
    wire [131:0] _1331;
    wire [63:0] _1332;
    wire [63:0] _1387;
    wire [63:0] data_75;
    wire [63:0] data_76;
    wire [63:0] data_77;
    wire [63:0] data_78;
    wire [5:0] address_80;
    wire _1312;
    wire read_enable_66;
    wire _1309;
    wire _1310;
    wire write_enable_80;
    wire _1314;
    wire [5:0] address_81;
    wire _1305;
    wire read_enable_67;
    wire _1302;
    wire _1303;
    wire write_enable_81;
    wire _1307;
    wire [131:0] _1317;
    wire [63:0] _1318;
    wire _1300 = 1'b0;
    wire _1299 = 1'b0;
    wire _1388;
    wire _53;
    reg PHASE_18;
    wire [63:0] q0_5;
    wire _1297 = 1'b0;
    wire _1296 = 1'b0;
    reg _1298;
    wire [63:0] _1377;
    wire [191:0] _1386;
    wire [63:0] _1389;
    wire [63:0] data_79;
    wire [63:0] data_80;
    wire [63:0] data_81;
    wire [63:0] data_82;
    wire [5:0] address_82;
    wire _1453;
    wire _1452;
    wire read_enable_68;
    wire _1446 = 1'b0;
    wire _1445 = 1'b0;
    wire _1443 = 1'b0;
    wire _1442 = 1'b0;
    wire _1440 = 1'b0;
    wire _1439 = 1'b0;
    wire _1437 = 1'b0;
    wire _1436 = 1'b0;
    wire _1434 = 1'b0;
    wire _1433 = 1'b0;
    wire _1431 = 1'b0;
    wire _1430 = 1'b0;
    wire _1428 = 1'b0;
    wire _1427 = 1'b0;
    wire _1425 = 1'b0;
    wire _1424 = 1'b0;
    wire _1422 = 1'b0;
    wire _1421 = 1'b0;
    reg _1423;
    reg _1426;
    reg _1429;
    reg _1432;
    reg _1435;
    reg _1438;
    reg _1441;
    reg _1444;
    reg _1447;
    wire _1448;
    wire _1419 = 1'b0;
    wire _1418 = 1'b0;
    wire _1416 = 1'b0;
    wire _1415 = 1'b0;
    wire _1413 = 1'b0;
    wire _1412 = 1'b0;
    wire _1410 = 1'b0;
    wire _1409 = 1'b0;
    wire _1407 = 1'b0;
    wire _1406 = 1'b0;
    wire _1404 = 1'b0;
    wire _1403 = 1'b0;
    wire _1401 = 1'b0;
    wire _1400 = 1'b0;
    wire _1398 = 1'b0;
    wire _1397 = 1'b0;
    wire _1395 = 1'b0;
    wire _1394 = 1'b0;
    reg _1396;
    reg _1399;
    reg _1402;
    reg _1405;
    reg _1408;
    reg _1411;
    reg _1414;
    reg _1417;
    reg _1420;
    wire _1449;
    wire _1450;
    wire write_enable_82;
    wire _1455;
    wire [131:0] _1462;
    wire [63:0] _1463;
    wire _1391 = 1'b0;
    wire _1390 = 1'b0;
    wire _1393;
    wire _55;
    reg PHASE_19;
    wire [63:0] _1475;
    wire [5:0] address_83;
    wire write_enable_83;
    wire [5:0] address_84;
    wire _1650;
    wire read_enable_69;
    wire _1648;
    wire write_enable_84;
    wire _1652;
    wire [131:0] _1657;
    wire [63:0] _1658;
    wire [5:0] _1643 = 6'b000000;
    wire [5:0] address_85;
    wire _1641;
    wire write_enable_85;
    wire [3:0] _280;
    wire _279;
    wire _277;
    wire [63:0] _276;
    wire [63:0] _275;
    wire [63:0] _274;
    wire [63:0] _273;
    wire [63:0] _272;
    wire [63:0] _271;
    wire [63:0] _270;
    wire [63:0] _1566;
    wire [63:0] _1565;
    wire [63:0] _1567;
    wire [63:0] _1563;
    wire [63:0] _1562;
    wire [63:0] q1_6;
    wire [63:0] _1568;
    wire [5:0] address_86;
    wire write_enable_86 = 1'b0;
    wire _1553;
    wire read_enable_70;
    wire [5:0] address_87;
    wire _1549;
    wire read_enable_71;
    wire _1547;
    wire write_enable_87;
    wire _1551;
    wire [131:0] _1558;
    wire [63:0] _1559;
    wire [63:0] data_83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_84;
    wire [5:0] _1541 = 6'b000000;
    wire _1539;
    wire _1538;
    wire _1537;
    wire _1536;
    wire _1535;
    wire _1534;
    wire [5:0] _1540;
    wire [5:0] address_88;
    wire write_enable_88 = 1'b0;
    wire _1531;
    wire read_enable_72;
    wire [63:0] data_85;
    wire [63:0] data_86;
    wire [5:0] _60;
    wire _1528;
    wire _1527;
    wire _1526;
    wire _1525;
    wire _1524;
    wire _1523;
    wire [5:0] _1529;
    wire [5:0] address_89;
    wire _1520;
    wire read_enable_73;
    wire [7:0] _62;
    wire _1518;
    wire write_enable_89;
    wire _1522;
    wire [131:0] _1545;
    wire [63:0] _1546;
    wire _1477 = 1'b0;
    wire _1476 = 1'b0;
    wire _1479;
    wire _63;
    reg PHASE_20;
    wire [63:0] _1560;
    wire [5:0] address_90;
    wire _1510;
    wire read_enable_74;
    wire write_enable_90;
    wire _1512;
    wire [5:0] address_91;
    wire _1505;
    wire read_enable_75;
    wire _1503;
    wire write_enable_91;
    wire _1507;
    wire [131:0] _1515;
    wire [63:0] _1516;
    wire [63:0] _1571;
    wire [63:0] data_87;
    wire [63:0] data_88;
    wire [63:0] data_89;
    wire [63:0] data_90;
    wire [5:0] _198 = 6'b000000;
    wire [5:0] _197 = 6'b000000;
    wire [5:0] _195 = 6'b000000;
    wire [5:0] _194 = 6'b000000;
    wire [5:0] _192 = 6'b000000;
    wire [5:0] _191 = 6'b000000;
    wire [5:0] _189 = 6'b000000;
    wire [5:0] _188 = 6'b000000;
    wire [5:0] _186 = 6'b000000;
    wire [5:0] _185 = 6'b000000;
    wire [5:0] _183 = 6'b000000;
    wire [5:0] _182 = 6'b000000;
    wire [5:0] _180 = 6'b000000;
    wire [5:0] _179 = 6'b000000;
    wire [5:0] _177 = 6'b000000;
    wire [5:0] _176 = 6'b000000;
    wire [5:0] _174 = 6'b000000;
    wire [5:0] _173 = 6'b000000;
    reg [5:0] _175;
    reg [5:0] _178;
    reg [5:0] _181;
    reg [5:0] _184;
    reg [5:0] _187;
    reg [5:0] _190;
    reg [5:0] _193;
    reg [5:0] _196;
    reg [5:0] _199;
    wire [5:0] _172;
    wire [5:0] address_92;
    wire _1496;
    wire read_enable_76;
    wire _1493;
    wire _1494;
    wire write_enable_92;
    wire _1498;
    wire [5:0] address_93;
    wire _1489;
    wire read_enable_77;
    wire _1486;
    wire _1487;
    wire write_enable_93;
    wire _1491;
    wire [131:0] _1501;
    wire [63:0] _1502;
    wire _99;
    wire _1484 = 1'b0;
    wire _1483 = 1'b0;
    wire _1572;
    wire _65;
    reg PHASE_21;
    wire [63:0] q0_6;
    wire _1481 = 1'b0;
    wire _1480 = 1'b0;
    wire _92;
    reg _1482;
    wire [63:0] _1561;
    wire [191:0] _1570;
    wire [63:0] _1573;
    wire [63:0] data_91;
    wire [63:0] data_92;
    wire [63:0] data_93;
    wire [63:0] data_94;
    wire [5:0] _163 = 6'b000000;
    wire [5:0] _162 = 6'b000000;
    wire [5:0] _160 = 6'b000000;
    wire [5:0] _159 = 6'b000000;
    wire [5:0] _157 = 6'b000000;
    wire [5:0] _156 = 6'b000000;
    wire [5:0] _154 = 6'b000000;
    wire [5:0] _153 = 6'b000000;
    wire [5:0] _151 = 6'b000000;
    wire [5:0] _150 = 6'b000000;
    wire [5:0] _148 = 6'b000000;
    wire [5:0] _147 = 6'b000000;
    wire [5:0] _145 = 6'b000000;
    wire [5:0] _144 = 6'b000000;
    wire [5:0] _142 = 6'b000000;
    wire [5:0] _141 = 6'b000000;
    wire [5:0] _139 = 6'b000000;
    wire [5:0] _138 = 6'b000000;
    wire [5:0] _137;
    reg [5:0] _140;
    reg [5:0] _143;
    reg [5:0] _146;
    reg [5:0] _149;
    reg [5:0] _152;
    reg [5:0] _155;
    reg [5:0] _158;
    reg [5:0] _161;
    reg [5:0] _164;
    wire [5:0] _68;
    wire [5:0] address_94;
    wire _1637;
    wire [7:0] _70;
    wire _1636;
    wire read_enable_78;
    wire _1630 = 1'b0;
    wire _1629 = 1'b0;
    wire _1627 = 1'b0;
    wire _1626 = 1'b0;
    wire _1624 = 1'b0;
    wire _1623 = 1'b0;
    wire _1621 = 1'b0;
    wire _1620 = 1'b0;
    wire _1618 = 1'b0;
    wire _1617 = 1'b0;
    wire _1615 = 1'b0;
    wire _1614 = 1'b0;
    wire _1612 = 1'b0;
    wire _1611 = 1'b0;
    wire _1609 = 1'b0;
    wire _1608 = 1'b0;
    wire _1606 = 1'b0;
    wire _1605 = 1'b0;
    wire _278;
    reg _1607;
    reg _1610;
    reg _1613;
    reg _1616;
    reg _1619;
    reg _1622;
    reg _1625;
    reg _1628;
    reg _1631;
    wire _1632;
    wire _1603 = 1'b0;
    wire _1602 = 1'b0;
    wire _1600 = 1'b0;
    wire _1599 = 1'b0;
    wire _1597 = 1'b0;
    wire _1596 = 1'b0;
    wire _1594 = 1'b0;
    wire _1593 = 1'b0;
    wire _1591 = 1'b0;
    wire _1590 = 1'b0;
    wire _1588 = 1'b0;
    wire _1587 = 1'b0;
    wire _1585 = 1'b0;
    wire _1584 = 1'b0;
    wire _1582 = 1'b0;
    wire _1581 = 1'b0;
    wire _1579 = 1'b0;
    wire _1578 = 1'b0;
    wire _130;
    reg _1580;
    reg _1583;
    reg _1586;
    reg _1589;
    reg _1592;
    reg _1595;
    reg _1598;
    reg _1601;
    reg _1604;
    wire _1633;
    wire _128 = 1'b0;
    wire _127 = 1'b0;
    wire _125 = 1'b0;
    wire _124 = 1'b0;
    wire _122 = 1'b0;
    wire _121 = 1'b0;
    wire _119 = 1'b0;
    wire _118 = 1'b0;
    wire _116 = 1'b0;
    wire _115 = 1'b0;
    wire _113 = 1'b0;
    wire _112 = 1'b0;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire vdd = 1'b1;
    wire _104 = 1'b0;
    wire _103 = 1'b0;
    wire _102;
    reg _105;
    reg _108;
    reg _111;
    reg _114;
    reg _117;
    reg _120;
    reg _123;
    reg _126;
    reg _129;
    wire _1634;
    wire write_enable_94;
    wire _1639;
    wire gnd = 1'b0;
    wire [131:0] _1646;
    wire [63:0] _1647;
    wire _72;
    wire _1575 = 1'b0;
    wire _1574 = 1'b0;
    wire _1577;
    wire _73;
    reg PHASE_22;
    wire [63:0] _1659;
    wire _76;
    wire _78;
    wire _80;
    wire _82;
    wire _84;
    wire [492:0] _91;
    wire _1660;

    /* logic */
    assign address = _360 ? _199 : _355;
    assign write_enable = _353 & _360;
    assign address_0 = _360 ? _164 : _68;
    assign _362 = ~ _360;
    assign read_enable = _348 & _362;
    assign _360 = ~ PHASE_1;
    assign write_enable_0 = _346 & _360;
    assign _364 = write_enable_0 | read_enable;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_364), .regcea(vdd), .wea(write_enable_0), .addra(address_0), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable), .regceb(vdd), .web(write_enable), .addrb(address), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_369[131:131]), .sbiterrb(_369[130:130]), .doutb(_369[129:66]), .dbiterra(_369[65:65]), .sbiterra(_369[64:64]), .douta(_369[63:0]) );
    assign _370 = _369[63:0];
    assign address_1 = PHASE_1 ? _199 : _355;
    assign _353 = _129 & _316;
    assign write_enable_1 = _353 & PHASE_1;
    assign _267 = _259[129:66];
    assign _266 = _246[129:66];
    assign _268 = PHASE ? _267 : _266;
    assign _264 = _216[129:66];
    assign _263 = _202[129:66];
    assign q1 = PHASE_0 ? _264 : _263;
    assign _269 = _96 ? _268 : q1;
    assign address_2 = _248 ? _242 : _241;
    assign _254 = ~ _248;
    assign read_enable_0 = _102 & _254;
    assign address_3 = _248 ? _60 : _230;
    assign _250 = ~ _248;
    assign read_enable_1 = _102 & _250;
    assign _248 = ~ PHASE;
    assign write_enable_3 = _219 & _248;
    assign _252 = write_enable_3 | read_enable_1;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_0
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_252), .regcea(vdd), .wea(write_enable_3), .addra(address_3), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_0), .regceb(vdd), .web(write_enable_2), .addrb(address_2), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_259[131:131]), .sbiterrb(_259[130:130]), .doutb(_259[129:66]), .dbiterra(_259[65:65]), .sbiterra(_259[64:64]), .douta(_259[63:0]) );
    assign _260 = _259[63:0];
    assign _240 = _172[5:5];
    assign _239 = _172[4:4];
    assign _238 = _172[3:3];
    assign _237 = _172[2:2];
    assign _236 = _172[1:1];
    assign _235 = _172[0:0];
    assign _241 = { _235, _236, _237, _238, _239, _240 };
    assign address_4 = PHASE ? _242 : _241;
    assign _232 = ~ PHASE;
    assign read_enable_2 = _102 & _232;
    assign data_1 = wr_d7;
    assign _229 = _137[5:5];
    assign _228 = _137[4:4];
    assign _227 = _137[3:3];
    assign _226 = _137[2:2];
    assign _225 = _137[1:1];
    assign _224 = _137[0:0];
    assign _230 = { _224, _225, _226, _227, _228, _229 };
    assign address_5 = PHASE ? _60 : _230;
    assign _221 = ~ PHASE;
    assign read_enable_3 = _102 & _221;
    assign _219 = _62[7:7];
    assign write_enable_5 = _219 & PHASE;
    assign _223 = write_enable_5 | read_enable_3;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_1
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_223), .regcea(vdd), .wea(write_enable_5), .addra(address_5), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_2), .regceb(vdd), .web(write_enable_4), .addrb(address_4), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_246[131:131]), .sbiterrb(_246[130:130]), .doutb(_246[129:66]), .dbiterra(_246[65:65]), .sbiterra(_246[64:64]), .douta(_246[63:0]) );
    assign _247 = _246[63:0];
    assign _89 = ~ PHASE;
    assign _3 = _89;
    always @(posedge _84) begin
        if (_82)
            PHASE <= _87;
        else
            if (_72)
                PHASE <= _3;
    end
    assign _261 = PHASE ? _260 : _247;
    assign address_6 = _204 ? _199 : _172;
    assign _211 = ~ _204;
    assign read_enable_4 = _102 & _211;
    assign write_enable_6 = _167 & _204;
    assign _213 = write_enable_6 | read_enable_4;
    assign address_7 = _204 ? _164 : _137;
    assign _206 = ~ _204;
    assign read_enable_5 = _102 & _206;
    assign _204 = ~ PHASE_0;
    assign write_enable_7 = _132 & _204;
    assign _208 = write_enable_7 | read_enable_5;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_2
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_208), .regcea(vdd), .wea(write_enable_7), .addra(address_7), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_213), .regceb(vdd), .web(write_enable_6), .addrb(address_6), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_216[131:131]), .sbiterrb(_216[130:130]), .doutb(_216[129:66]), .dbiterra(_216[65:65]), .sbiterra(_216[64:64]), .douta(_216[63:0]) );
    assign _217 = _216[63:0];
    assign _283 = _282[127:64];
    assign data_3 = _283;
    assign address_8 = PHASE_0 ? _199 : _172;
    assign _169 = ~ PHASE_0;
    assign read_enable_6 = _102 & _169;
    assign _166 = ~ _130;
    assign _167 = _129 & _166;
    assign write_enable_8 = _167 & PHASE_0;
    assign _171 = write_enable_8 | read_enable_6;
    assign address_9 = PHASE_0 ? _164 : _137;
    assign _134 = ~ PHASE_0;
    assign read_enable_7 = _102 & _134;
    assign _131 = ~ _130;
    assign _132 = _129 & _131;
    assign write_enable_9 = _132 & PHASE_0;
    assign _136 = write_enable_9 | read_enable_7;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_3
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_136), .regcea(vdd), .wea(write_enable_9), .addra(address_9), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_171), .regceb(vdd), .web(write_enable_8), .addrb(address_8), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_202[131:131]), .sbiterrb(_202[130:130]), .doutb(_202[129:66]), .dbiterra(_202[65:65]), .sbiterra(_202[64:64]), .douta(_202[63:0]) );
    assign _203 = _202[63:0];
    assign _284 = ~ PHASE_0;
    assign _5 = _284;
    always @(posedge _84) begin
        if (_82)
            PHASE_0 <= _98;
        else
            if (_99)
                PHASE_0 <= _5;
    end
    assign q0 = PHASE_0 ? _217 : _203;
    always @(posedge _84) begin
        if (_82)
            _96 <= _94;
        else
            _96 <= _92;
    end
    assign _262 = _96 ? _261 : q0;
    dp_30
        dp_6
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_262), .d2(_269), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_282[191:128]), .q2(_282[127:64]), .q1(_282[63:0]) );
    assign _285 = _282[63:0];
    assign data_7 = _285;
    assign address_10 = PHASE_1 ? _164 : _68;
    assign _349 = ~ PHASE_1;
    assign _348 = _70[7:7];
    assign read_enable_8 = _348 & _349;
    always @(posedge _84) begin
        if (_82)
            _319 <= _318;
        else
            _319 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _322 <= _321;
        else
            _322 <= _319;
    end
    always @(posedge _84) begin
        if (_82)
            _325 <= _324;
        else
            _325 <= _322;
    end
    always @(posedge _84) begin
        if (_82)
            _328 <= _327;
        else
            _328 <= _325;
    end
    always @(posedge _84) begin
        if (_82)
            _331 <= _330;
        else
            _331 <= _328;
    end
    always @(posedge _84) begin
        if (_82)
            _334 <= _333;
        else
            _334 <= _331;
    end
    always @(posedge _84) begin
        if (_82)
            _337 <= _336;
        else
            _337 <= _334;
    end
    always @(posedge _84) begin
        if (_82)
            _340 <= _339;
        else
            _340 <= _337;
    end
    always @(posedge _84) begin
        if (_82)
            _343 <= _342;
        else
            _343 <= _340;
    end
    assign _344 = ~ _343;
    always @(posedge _84) begin
        if (_82)
            _292 <= _291;
        else
            _292 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _295 <= _294;
        else
            _295 <= _292;
    end
    always @(posedge _84) begin
        if (_82)
            _298 <= _297;
        else
            _298 <= _295;
    end
    always @(posedge _84) begin
        if (_82)
            _301 <= _300;
        else
            _301 <= _298;
    end
    always @(posedge _84) begin
        if (_82)
            _304 <= _303;
        else
            _304 <= _301;
    end
    always @(posedge _84) begin
        if (_82)
            _307 <= _306;
        else
            _307 <= _304;
    end
    always @(posedge _84) begin
        if (_82)
            _310 <= _309;
        else
            _310 <= _307;
    end
    always @(posedge _84) begin
        if (_82)
            _313 <= _312;
        else
            _313 <= _310;
    end
    always @(posedge _84) begin
        if (_82)
            _316 <= _315;
        else
            _316 <= _313;
    end
    assign _345 = _316 & _344;
    assign _346 = _129 & _345;
    assign write_enable_10 = _346 & PHASE_1;
    assign _351 = write_enable_10 | read_enable_8;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_4
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_351), .regcea(vdd), .wea(write_enable_10), .addra(address_10), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_1), .regceb(vdd), .web(write_enable_1), .addrb(address_1), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_358[131:131]), .sbiterrb(_358[130:130]), .doutb(_358[129:66]), .dbiterra(_358[65:65]), .sbiterra(_358[64:64]), .douta(_358[63:0]) );
    assign _359 = _358[63:0];
    assign _289 = ~ PHASE_1;
    assign _7 = _289;
    always @(posedge _84) begin
        if (_82)
            PHASE_1 <= _287;
        else
            if (_72)
                PHASE_1 <= _7;
    end
    assign _371 = PHASE_1 ? _370 : _359;
    assign address_11 = _544 ? _199 : _539;
    assign write_enable_11 = _537 & _544;
    assign address_12 = _544 ? _164 : _68;
    assign _546 = ~ _544;
    assign read_enable_9 = _532 & _546;
    assign _544 = ~ PHASE_4;
    assign write_enable_12 = _530 & _544;
    assign _548 = write_enable_12 | read_enable_9;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_5
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_548), .regcea(vdd), .wea(write_enable_12), .addra(address_12), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_11), .regceb(vdd), .web(write_enable_11), .addrb(address_11), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_553[131:131]), .sbiterrb(_553[130:130]), .doutb(_553[129:66]), .dbiterra(_553[65:65]), .sbiterra(_553[64:64]), .douta(_553[63:0]) );
    assign _554 = _553[63:0];
    assign address_13 = PHASE_4 ? _199 : _539;
    assign _537 = _129 & _500;
    assign write_enable_13 = _537 & PHASE_4;
    assign _462 = _454[129:66];
    assign _461 = _441[129:66];
    assign _463 = PHASE_2 ? _462 : _461;
    assign _459 = _411[129:66];
    assign _458 = _397[129:66];
    assign q1_0 = PHASE_3 ? _459 : _458;
    assign _464 = _378 ? _463 : q1_0;
    assign address_14 = _443 ? _437 : _436;
    assign _449 = ~ _443;
    assign read_enable_10 = _102 & _449;
    assign address_15 = _443 ? _60 : _425;
    assign _445 = ~ _443;
    assign read_enable_11 = _102 & _445;
    assign _443 = ~ PHASE_2;
    assign write_enable_15 = _414 & _443;
    assign _447 = write_enable_15 | read_enable_11;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_6
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_447), .regcea(vdd), .wea(write_enable_15), .addra(address_15), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_10), .regceb(vdd), .web(write_enable_14), .addrb(address_14), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_454[131:131]), .sbiterrb(_454[130:130]), .doutb(_454[129:66]), .dbiterra(_454[65:65]), .sbiterra(_454[64:64]), .douta(_454[63:0]) );
    assign _455 = _454[63:0];
    assign _435 = _172[5:5];
    assign _434 = _172[4:4];
    assign _433 = _172[3:3];
    assign _432 = _172[2:2];
    assign _431 = _172[1:1];
    assign _430 = _172[0:0];
    assign _436 = { _430, _431, _432, _433, _434, _435 };
    assign address_16 = PHASE_2 ? _437 : _436;
    assign _427 = ~ PHASE_2;
    assign read_enable_12 = _102 & _427;
    assign data_13 = wr_d6;
    assign _424 = _137[5:5];
    assign _423 = _137[4:4];
    assign _422 = _137[3:3];
    assign _421 = _137[2:2];
    assign _420 = _137[1:1];
    assign _419 = _137[0:0];
    assign _425 = { _419, _420, _421, _422, _423, _424 };
    assign address_17 = PHASE_2 ? _60 : _425;
    assign _416 = ~ PHASE_2;
    assign read_enable_13 = _102 & _416;
    assign _414 = _62[6:6];
    assign write_enable_17 = _414 & PHASE_2;
    assign _418 = write_enable_17 | read_enable_13;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_7
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_418), .regcea(vdd), .wea(write_enable_17), .addra(address_17), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_12), .regceb(vdd), .web(write_enable_16), .addrb(address_16), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_441[131:131]), .sbiterrb(_441[130:130]), .doutb(_441[129:66]), .dbiterra(_441[65:65]), .sbiterra(_441[64:64]), .douta(_441[63:0]) );
    assign _442 = _441[63:0];
    assign _375 = ~ PHASE_2;
    assign _11 = _375;
    always @(posedge _84) begin
        if (_82)
            PHASE_2 <= _373;
        else
            if (_72)
                PHASE_2 <= _11;
    end
    assign _456 = PHASE_2 ? _455 : _442;
    assign address_18 = _399 ? _199 : _172;
    assign _406 = ~ _399;
    assign read_enable_14 = _102 & _406;
    assign write_enable_18 = _390 & _399;
    assign _408 = write_enable_18 | read_enable_14;
    assign address_19 = _399 ? _164 : _137;
    assign _401 = ~ _399;
    assign read_enable_15 = _102 & _401;
    assign _399 = ~ PHASE_3;
    assign write_enable_19 = _383 & _399;
    assign _403 = write_enable_19 | read_enable_15;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_8
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_403), .regcea(vdd), .wea(write_enable_19), .addra(address_19), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_408), .regceb(vdd), .web(write_enable_18), .addrb(address_18), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_411[131:131]), .sbiterrb(_411[130:130]), .doutb(_411[129:66]), .dbiterra(_411[65:65]), .sbiterra(_411[64:64]), .douta(_411[63:0]) );
    assign _412 = _411[63:0];
    assign _467 = _466[127:64];
    assign data_15 = _467;
    assign address_20 = PHASE_3 ? _199 : _172;
    assign _392 = ~ PHASE_3;
    assign read_enable_16 = _102 & _392;
    assign _389 = ~ _130;
    assign _390 = _129 & _389;
    assign write_enable_20 = _390 & PHASE_3;
    assign _394 = write_enable_20 | read_enable_16;
    assign address_21 = PHASE_3 ? _164 : _137;
    assign _385 = ~ PHASE_3;
    assign read_enable_17 = _102 & _385;
    assign _382 = ~ _130;
    assign _383 = _129 & _382;
    assign write_enable_21 = _383 & PHASE_3;
    assign _387 = write_enable_21 | read_enable_17;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_9
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_387), .regcea(vdd), .wea(write_enable_21), .addra(address_21), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_394), .regceb(vdd), .web(write_enable_20), .addrb(address_20), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_397[131:131]), .sbiterrb(_397[130:130]), .doutb(_397[129:66]), .dbiterra(_397[65:65]), .sbiterra(_397[64:64]), .douta(_397[63:0]) );
    assign _398 = _397[63:0];
    assign _468 = ~ PHASE_3;
    assign _13 = _468;
    always @(posedge _84) begin
        if (_82)
            PHASE_3 <= _380;
        else
            if (_99)
                PHASE_3 <= _13;
    end
    assign q0_0 = PHASE_3 ? _412 : _398;
    always @(posedge _84) begin
        if (_82)
            _378 <= _377;
        else
            _378 <= _92;
    end
    assign _457 = _378 ? _456 : q0_0;
    dp_29
        dp_5
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_457), .d2(_464), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_466[191:128]), .q2(_466[127:64]), .q1(_466[63:0]) );
    assign _469 = _466[63:0];
    assign data_19 = _469;
    assign address_22 = PHASE_4 ? _164 : _68;
    assign _533 = ~ PHASE_4;
    assign _532 = _70[6:6];
    assign read_enable_18 = _532 & _533;
    always @(posedge _84) begin
        if (_82)
            _503 <= _502;
        else
            _503 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _506 <= _505;
        else
            _506 <= _503;
    end
    always @(posedge _84) begin
        if (_82)
            _509 <= _508;
        else
            _509 <= _506;
    end
    always @(posedge _84) begin
        if (_82)
            _512 <= _511;
        else
            _512 <= _509;
    end
    always @(posedge _84) begin
        if (_82)
            _515 <= _514;
        else
            _515 <= _512;
    end
    always @(posedge _84) begin
        if (_82)
            _518 <= _517;
        else
            _518 <= _515;
    end
    always @(posedge _84) begin
        if (_82)
            _521 <= _520;
        else
            _521 <= _518;
    end
    always @(posedge _84) begin
        if (_82)
            _524 <= _523;
        else
            _524 <= _521;
    end
    always @(posedge _84) begin
        if (_82)
            _527 <= _526;
        else
            _527 <= _524;
    end
    assign _528 = ~ _527;
    always @(posedge _84) begin
        if (_82)
            _476 <= _475;
        else
            _476 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _479 <= _478;
        else
            _479 <= _476;
    end
    always @(posedge _84) begin
        if (_82)
            _482 <= _481;
        else
            _482 <= _479;
    end
    always @(posedge _84) begin
        if (_82)
            _485 <= _484;
        else
            _485 <= _482;
    end
    always @(posedge _84) begin
        if (_82)
            _488 <= _487;
        else
            _488 <= _485;
    end
    always @(posedge _84) begin
        if (_82)
            _491 <= _490;
        else
            _491 <= _488;
    end
    always @(posedge _84) begin
        if (_82)
            _494 <= _493;
        else
            _494 <= _491;
    end
    always @(posedge _84) begin
        if (_82)
            _497 <= _496;
        else
            _497 <= _494;
    end
    always @(posedge _84) begin
        if (_82)
            _500 <= _499;
        else
            _500 <= _497;
    end
    assign _529 = _500 & _528;
    assign _530 = _129 & _529;
    assign write_enable_22 = _530 & PHASE_4;
    assign _535 = write_enable_22 | read_enable_18;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_10
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_535), .regcea(vdd), .wea(write_enable_22), .addra(address_22), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_13), .regceb(vdd), .web(write_enable_13), .addrb(address_13), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_542[131:131]), .sbiterrb(_542[130:130]), .doutb(_542[129:66]), .dbiterra(_542[65:65]), .sbiterra(_542[64:64]), .douta(_542[63:0]) );
    assign _543 = _542[63:0];
    assign _473 = ~ PHASE_4;
    assign _15 = _473;
    always @(posedge _84) begin
        if (_82)
            PHASE_4 <= _471;
        else
            if (_72)
                PHASE_4 <= _15;
    end
    assign _555 = PHASE_4 ? _554 : _543;
    assign address_23 = _728 ? _199 : _723;
    assign write_enable_23 = _721 & _728;
    assign address_24 = _728 ? _164 : _68;
    assign _730 = ~ _728;
    assign read_enable_19 = _716 & _730;
    assign _728 = ~ PHASE_7;
    assign write_enable_24 = _714 & _728;
    assign _732 = write_enable_24 | read_enable_19;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_11
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_732), .regcea(vdd), .wea(write_enable_24), .addra(address_24), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_23), .regceb(vdd), .web(write_enable_23), .addrb(address_23), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_737[131:131]), .sbiterrb(_737[130:130]), .doutb(_737[129:66]), .dbiterra(_737[65:65]), .sbiterra(_737[64:64]), .douta(_737[63:0]) );
    assign _738 = _737[63:0];
    assign address_25 = PHASE_7 ? _199 : _723;
    assign _721 = _129 & _684;
    assign write_enable_25 = _721 & PHASE_7;
    assign _646 = _638[129:66];
    assign _645 = _625[129:66];
    assign _647 = PHASE_5 ? _646 : _645;
    assign _643 = _595[129:66];
    assign _642 = _581[129:66];
    assign q1_1 = PHASE_6 ? _643 : _642;
    assign _648 = _562 ? _647 : q1_1;
    assign address_26 = _627 ? _621 : _620;
    assign _633 = ~ _627;
    assign read_enable_20 = _102 & _633;
    assign address_27 = _627 ? _60 : _609;
    assign _629 = ~ _627;
    assign read_enable_21 = _102 & _629;
    assign _627 = ~ PHASE_5;
    assign write_enable_27 = _598 & _627;
    assign _631 = write_enable_27 | read_enable_21;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_12
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_631), .regcea(vdd), .wea(write_enable_27), .addra(address_27), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_20), .regceb(vdd), .web(write_enable_26), .addrb(address_26), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_638[131:131]), .sbiterrb(_638[130:130]), .doutb(_638[129:66]), .dbiterra(_638[65:65]), .sbiterra(_638[64:64]), .douta(_638[63:0]) );
    assign _639 = _638[63:0];
    assign _619 = _172[5:5];
    assign _618 = _172[4:4];
    assign _617 = _172[3:3];
    assign _616 = _172[2:2];
    assign _615 = _172[1:1];
    assign _614 = _172[0:0];
    assign _620 = { _614, _615, _616, _617, _618, _619 };
    assign address_28 = PHASE_5 ? _621 : _620;
    assign _611 = ~ PHASE_5;
    assign read_enable_22 = _102 & _611;
    assign data_25 = wr_d5;
    assign _608 = _137[5:5];
    assign _607 = _137[4:4];
    assign _606 = _137[3:3];
    assign _605 = _137[2:2];
    assign _604 = _137[1:1];
    assign _603 = _137[0:0];
    assign _609 = { _603, _604, _605, _606, _607, _608 };
    assign address_29 = PHASE_5 ? _60 : _609;
    assign _600 = ~ PHASE_5;
    assign read_enable_23 = _102 & _600;
    assign _598 = _62[5:5];
    assign write_enable_29 = _598 & PHASE_5;
    assign _602 = write_enable_29 | read_enable_23;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_13
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_602), .regcea(vdd), .wea(write_enable_29), .addra(address_29), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_22), .regceb(vdd), .web(write_enable_28), .addrb(address_28), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_625[131:131]), .sbiterrb(_625[130:130]), .doutb(_625[129:66]), .dbiterra(_625[65:65]), .sbiterra(_625[64:64]), .douta(_625[63:0]) );
    assign _626 = _625[63:0];
    assign _559 = ~ PHASE_5;
    assign _19 = _559;
    always @(posedge _84) begin
        if (_82)
            PHASE_5 <= _557;
        else
            if (_72)
                PHASE_5 <= _19;
    end
    assign _640 = PHASE_5 ? _639 : _626;
    assign address_30 = _583 ? _199 : _172;
    assign _590 = ~ _583;
    assign read_enable_24 = _102 & _590;
    assign write_enable_30 = _574 & _583;
    assign _592 = write_enable_30 | read_enable_24;
    assign address_31 = _583 ? _164 : _137;
    assign _585 = ~ _583;
    assign read_enable_25 = _102 & _585;
    assign _583 = ~ PHASE_6;
    assign write_enable_31 = _567 & _583;
    assign _587 = write_enable_31 | read_enable_25;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_14
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_587), .regcea(vdd), .wea(write_enable_31), .addra(address_31), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_592), .regceb(vdd), .web(write_enable_30), .addrb(address_30), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_595[131:131]), .sbiterrb(_595[130:130]), .doutb(_595[129:66]), .dbiterra(_595[65:65]), .sbiterra(_595[64:64]), .douta(_595[63:0]) );
    assign _596 = _595[63:0];
    assign _651 = _650[127:64];
    assign data_27 = _651;
    assign address_32 = PHASE_6 ? _199 : _172;
    assign _576 = ~ PHASE_6;
    assign read_enable_26 = _102 & _576;
    assign _573 = ~ _130;
    assign _574 = _129 & _573;
    assign write_enable_32 = _574 & PHASE_6;
    assign _578 = write_enable_32 | read_enable_26;
    assign address_33 = PHASE_6 ? _164 : _137;
    assign _569 = ~ PHASE_6;
    assign read_enable_27 = _102 & _569;
    assign _566 = ~ _130;
    assign _567 = _129 & _566;
    assign write_enable_33 = _567 & PHASE_6;
    assign _571 = write_enable_33 | read_enable_27;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_15
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_571), .regcea(vdd), .wea(write_enable_33), .addra(address_33), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_578), .regceb(vdd), .web(write_enable_32), .addrb(address_32), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_581[131:131]), .sbiterrb(_581[130:130]), .doutb(_581[129:66]), .dbiterra(_581[65:65]), .sbiterra(_581[64:64]), .douta(_581[63:0]) );
    assign _582 = _581[63:0];
    assign _652 = ~ PHASE_6;
    assign _21 = _652;
    always @(posedge _84) begin
        if (_82)
            PHASE_6 <= _564;
        else
            if (_99)
                PHASE_6 <= _21;
    end
    assign q0_1 = PHASE_6 ? _596 : _582;
    always @(posedge _84) begin
        if (_82)
            _562 <= _561;
        else
            _562 <= _92;
    end
    assign _641 = _562 ? _640 : q0_1;
    dp_28
        dp_4
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_641), .d2(_648), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_650[191:128]), .q2(_650[127:64]), .q1(_650[63:0]) );
    assign _653 = _650[63:0];
    assign data_31 = _653;
    assign address_34 = PHASE_7 ? _164 : _68;
    assign _717 = ~ PHASE_7;
    assign _716 = _70[5:5];
    assign read_enable_28 = _716 & _717;
    always @(posedge _84) begin
        if (_82)
            _687 <= _686;
        else
            _687 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _690 <= _689;
        else
            _690 <= _687;
    end
    always @(posedge _84) begin
        if (_82)
            _693 <= _692;
        else
            _693 <= _690;
    end
    always @(posedge _84) begin
        if (_82)
            _696 <= _695;
        else
            _696 <= _693;
    end
    always @(posedge _84) begin
        if (_82)
            _699 <= _698;
        else
            _699 <= _696;
    end
    always @(posedge _84) begin
        if (_82)
            _702 <= _701;
        else
            _702 <= _699;
    end
    always @(posedge _84) begin
        if (_82)
            _705 <= _704;
        else
            _705 <= _702;
    end
    always @(posedge _84) begin
        if (_82)
            _708 <= _707;
        else
            _708 <= _705;
    end
    always @(posedge _84) begin
        if (_82)
            _711 <= _710;
        else
            _711 <= _708;
    end
    assign _712 = ~ _711;
    always @(posedge _84) begin
        if (_82)
            _660 <= _659;
        else
            _660 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _663 <= _662;
        else
            _663 <= _660;
    end
    always @(posedge _84) begin
        if (_82)
            _666 <= _665;
        else
            _666 <= _663;
    end
    always @(posedge _84) begin
        if (_82)
            _669 <= _668;
        else
            _669 <= _666;
    end
    always @(posedge _84) begin
        if (_82)
            _672 <= _671;
        else
            _672 <= _669;
    end
    always @(posedge _84) begin
        if (_82)
            _675 <= _674;
        else
            _675 <= _672;
    end
    always @(posedge _84) begin
        if (_82)
            _678 <= _677;
        else
            _678 <= _675;
    end
    always @(posedge _84) begin
        if (_82)
            _681 <= _680;
        else
            _681 <= _678;
    end
    always @(posedge _84) begin
        if (_82)
            _684 <= _683;
        else
            _684 <= _681;
    end
    assign _713 = _684 & _712;
    assign _714 = _129 & _713;
    assign write_enable_34 = _714 & PHASE_7;
    assign _719 = write_enable_34 | read_enable_28;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_16
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_719), .regcea(vdd), .wea(write_enable_34), .addra(address_34), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_25), .regceb(vdd), .web(write_enable_25), .addrb(address_25), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_726[131:131]), .sbiterrb(_726[130:130]), .doutb(_726[129:66]), .dbiterra(_726[65:65]), .sbiterra(_726[64:64]), .douta(_726[63:0]) );
    assign _727 = _726[63:0];
    assign _657 = ~ PHASE_7;
    assign _23 = _657;
    always @(posedge _84) begin
        if (_82)
            PHASE_7 <= _655;
        else
            if (_72)
                PHASE_7 <= _23;
    end
    assign _739 = PHASE_7 ? _738 : _727;
    assign address_35 = _912 ? _199 : _907;
    assign write_enable_35 = _905 & _912;
    assign address_36 = _912 ? _164 : _68;
    assign _914 = ~ _912;
    assign read_enable_29 = _900 & _914;
    assign _912 = ~ PHASE_10;
    assign write_enable_36 = _898 & _912;
    assign _916 = write_enable_36 | read_enable_29;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_17
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_916), .regcea(vdd), .wea(write_enable_36), .addra(address_36), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_35), .regceb(vdd), .web(write_enable_35), .addrb(address_35), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_921[131:131]), .sbiterrb(_921[130:130]), .doutb(_921[129:66]), .dbiterra(_921[65:65]), .sbiterra(_921[64:64]), .douta(_921[63:0]) );
    assign _922 = _921[63:0];
    assign address_37 = PHASE_10 ? _199 : _907;
    assign _905 = _129 & _868;
    assign write_enable_37 = _905 & PHASE_10;
    assign _830 = _822[129:66];
    assign _829 = _809[129:66];
    assign _831 = PHASE_8 ? _830 : _829;
    assign _827 = _779[129:66];
    assign _826 = _765[129:66];
    assign q1_2 = PHASE_9 ? _827 : _826;
    assign _832 = _746 ? _831 : q1_2;
    assign address_38 = _811 ? _805 : _804;
    assign _817 = ~ _811;
    assign read_enable_30 = _102 & _817;
    assign address_39 = _811 ? _60 : _793;
    assign _813 = ~ _811;
    assign read_enable_31 = _102 & _813;
    assign _811 = ~ PHASE_8;
    assign write_enable_39 = _782 & _811;
    assign _815 = write_enable_39 | read_enable_31;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_18
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_815), .regcea(vdd), .wea(write_enable_39), .addra(address_39), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_30), .regceb(vdd), .web(write_enable_38), .addrb(address_38), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_822[131:131]), .sbiterrb(_822[130:130]), .doutb(_822[129:66]), .dbiterra(_822[65:65]), .sbiterra(_822[64:64]), .douta(_822[63:0]) );
    assign _823 = _822[63:0];
    assign _803 = _172[5:5];
    assign _802 = _172[4:4];
    assign _801 = _172[3:3];
    assign _800 = _172[2:2];
    assign _799 = _172[1:1];
    assign _798 = _172[0:0];
    assign _804 = { _798, _799, _800, _801, _802, _803 };
    assign address_40 = PHASE_8 ? _805 : _804;
    assign _795 = ~ PHASE_8;
    assign read_enable_32 = _102 & _795;
    assign data_37 = wr_d4;
    assign _792 = _137[5:5];
    assign _791 = _137[4:4];
    assign _790 = _137[3:3];
    assign _789 = _137[2:2];
    assign _788 = _137[1:1];
    assign _787 = _137[0:0];
    assign _793 = { _787, _788, _789, _790, _791, _792 };
    assign address_41 = PHASE_8 ? _60 : _793;
    assign _784 = ~ PHASE_8;
    assign read_enable_33 = _102 & _784;
    assign _782 = _62[4:4];
    assign write_enable_41 = _782 & PHASE_8;
    assign _786 = write_enable_41 | read_enable_33;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_19
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_786), .regcea(vdd), .wea(write_enable_41), .addra(address_41), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_32), .regceb(vdd), .web(write_enable_40), .addrb(address_40), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_809[131:131]), .sbiterrb(_809[130:130]), .doutb(_809[129:66]), .dbiterra(_809[65:65]), .sbiterra(_809[64:64]), .douta(_809[63:0]) );
    assign _810 = _809[63:0];
    assign _743 = ~ PHASE_8;
    assign _27 = _743;
    always @(posedge _84) begin
        if (_82)
            PHASE_8 <= _741;
        else
            if (_72)
                PHASE_8 <= _27;
    end
    assign _824 = PHASE_8 ? _823 : _810;
    assign address_42 = _767 ? _199 : _172;
    assign _774 = ~ _767;
    assign read_enable_34 = _102 & _774;
    assign write_enable_42 = _758 & _767;
    assign _776 = write_enable_42 | read_enable_34;
    assign address_43 = _767 ? _164 : _137;
    assign _769 = ~ _767;
    assign read_enable_35 = _102 & _769;
    assign _767 = ~ PHASE_9;
    assign write_enable_43 = _751 & _767;
    assign _771 = write_enable_43 | read_enable_35;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_20
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_771), .regcea(vdd), .wea(write_enable_43), .addra(address_43), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_776), .regceb(vdd), .web(write_enable_42), .addrb(address_42), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_779[131:131]), .sbiterrb(_779[130:130]), .doutb(_779[129:66]), .dbiterra(_779[65:65]), .sbiterra(_779[64:64]), .douta(_779[63:0]) );
    assign _780 = _779[63:0];
    assign _835 = _834[127:64];
    assign data_39 = _835;
    assign address_44 = PHASE_9 ? _199 : _172;
    assign _760 = ~ PHASE_9;
    assign read_enable_36 = _102 & _760;
    assign _757 = ~ _130;
    assign _758 = _129 & _757;
    assign write_enable_44 = _758 & PHASE_9;
    assign _762 = write_enable_44 | read_enable_36;
    assign address_45 = PHASE_9 ? _164 : _137;
    assign _753 = ~ PHASE_9;
    assign read_enable_37 = _102 & _753;
    assign _750 = ~ _130;
    assign _751 = _129 & _750;
    assign write_enable_45 = _751 & PHASE_9;
    assign _755 = write_enable_45 | read_enable_37;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_21
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_755), .regcea(vdd), .wea(write_enable_45), .addra(address_45), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_762), .regceb(vdd), .web(write_enable_44), .addrb(address_44), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_765[131:131]), .sbiterrb(_765[130:130]), .doutb(_765[129:66]), .dbiterra(_765[65:65]), .sbiterra(_765[64:64]), .douta(_765[63:0]) );
    assign _766 = _765[63:0];
    assign _836 = ~ PHASE_9;
    assign _29 = _836;
    always @(posedge _84) begin
        if (_82)
            PHASE_9 <= _748;
        else
            if (_99)
                PHASE_9 <= _29;
    end
    assign q0_2 = PHASE_9 ? _780 : _766;
    always @(posedge _84) begin
        if (_82)
            _746 <= _745;
        else
            _746 <= _92;
    end
    assign _825 = _746 ? _824 : q0_2;
    dp_27
        dp_3
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_825), .d2(_832), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_834[191:128]), .q2(_834[127:64]), .q1(_834[63:0]) );
    assign _837 = _834[63:0];
    assign data_43 = _837;
    assign address_46 = PHASE_10 ? _164 : _68;
    assign _901 = ~ PHASE_10;
    assign _900 = _70[4:4];
    assign read_enable_38 = _900 & _901;
    always @(posedge _84) begin
        if (_82)
            _871 <= _870;
        else
            _871 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _874 <= _873;
        else
            _874 <= _871;
    end
    always @(posedge _84) begin
        if (_82)
            _877 <= _876;
        else
            _877 <= _874;
    end
    always @(posedge _84) begin
        if (_82)
            _880 <= _879;
        else
            _880 <= _877;
    end
    always @(posedge _84) begin
        if (_82)
            _883 <= _882;
        else
            _883 <= _880;
    end
    always @(posedge _84) begin
        if (_82)
            _886 <= _885;
        else
            _886 <= _883;
    end
    always @(posedge _84) begin
        if (_82)
            _889 <= _888;
        else
            _889 <= _886;
    end
    always @(posedge _84) begin
        if (_82)
            _892 <= _891;
        else
            _892 <= _889;
    end
    always @(posedge _84) begin
        if (_82)
            _895 <= _894;
        else
            _895 <= _892;
    end
    assign _896 = ~ _895;
    always @(posedge _84) begin
        if (_82)
            _844 <= _843;
        else
            _844 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _847 <= _846;
        else
            _847 <= _844;
    end
    always @(posedge _84) begin
        if (_82)
            _850 <= _849;
        else
            _850 <= _847;
    end
    always @(posedge _84) begin
        if (_82)
            _853 <= _852;
        else
            _853 <= _850;
    end
    always @(posedge _84) begin
        if (_82)
            _856 <= _855;
        else
            _856 <= _853;
    end
    always @(posedge _84) begin
        if (_82)
            _859 <= _858;
        else
            _859 <= _856;
    end
    always @(posedge _84) begin
        if (_82)
            _862 <= _861;
        else
            _862 <= _859;
    end
    always @(posedge _84) begin
        if (_82)
            _865 <= _864;
        else
            _865 <= _862;
    end
    always @(posedge _84) begin
        if (_82)
            _868 <= _867;
        else
            _868 <= _865;
    end
    assign _897 = _868 & _896;
    assign _898 = _129 & _897;
    assign write_enable_46 = _898 & PHASE_10;
    assign _903 = write_enable_46 | read_enable_38;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_22
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_903), .regcea(vdd), .wea(write_enable_46), .addra(address_46), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_37), .regceb(vdd), .web(write_enable_37), .addrb(address_37), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_910[131:131]), .sbiterrb(_910[130:130]), .doutb(_910[129:66]), .dbiterra(_910[65:65]), .sbiterra(_910[64:64]), .douta(_910[63:0]) );
    assign _911 = _910[63:0];
    assign _841 = ~ PHASE_10;
    assign _31 = _841;
    always @(posedge _84) begin
        if (_82)
            PHASE_10 <= _839;
        else
            if (_72)
                PHASE_10 <= _31;
    end
    assign _923 = PHASE_10 ? _922 : _911;
    assign address_47 = _1096 ? _199 : _1091;
    assign write_enable_47 = _1089 & _1096;
    assign address_48 = _1096 ? _164 : _68;
    assign _1098 = ~ _1096;
    assign read_enable_39 = _1084 & _1098;
    assign _1096 = ~ PHASE_13;
    assign write_enable_48 = _1082 & _1096;
    assign _1100 = write_enable_48 | read_enable_39;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_23
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1100), .regcea(vdd), .wea(write_enable_48), .addra(address_48), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_47), .regceb(vdd), .web(write_enable_47), .addrb(address_47), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1105[131:131]), .sbiterrb(_1105[130:130]), .doutb(_1105[129:66]), .dbiterra(_1105[65:65]), .sbiterra(_1105[64:64]), .douta(_1105[63:0]) );
    assign _1106 = _1105[63:0];
    assign address_49 = PHASE_13 ? _199 : _1091;
    assign _1089 = _129 & _1052;
    assign write_enable_49 = _1089 & PHASE_13;
    assign _1014 = _1006[129:66];
    assign _1013 = _993[129:66];
    assign _1015 = PHASE_11 ? _1014 : _1013;
    assign _1011 = _963[129:66];
    assign _1010 = _949[129:66];
    assign q1_3 = PHASE_12 ? _1011 : _1010;
    assign _1016 = _930 ? _1015 : q1_3;
    assign address_50 = _995 ? _989 : _988;
    assign _1001 = ~ _995;
    assign read_enable_40 = _102 & _1001;
    assign address_51 = _995 ? _60 : _977;
    assign _997 = ~ _995;
    assign read_enable_41 = _102 & _997;
    assign _995 = ~ PHASE_11;
    assign write_enable_51 = _966 & _995;
    assign _999 = write_enable_51 | read_enable_41;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_24
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_999), .regcea(vdd), .wea(write_enable_51), .addra(address_51), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_40), .regceb(vdd), .web(write_enable_50), .addrb(address_50), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1006[131:131]), .sbiterrb(_1006[130:130]), .doutb(_1006[129:66]), .dbiterra(_1006[65:65]), .sbiterra(_1006[64:64]), .douta(_1006[63:0]) );
    assign _1007 = _1006[63:0];
    assign _987 = _172[5:5];
    assign _986 = _172[4:4];
    assign _985 = _172[3:3];
    assign _984 = _172[2:2];
    assign _983 = _172[1:1];
    assign _982 = _172[0:0];
    assign _988 = { _982, _983, _984, _985, _986, _987 };
    assign address_52 = PHASE_11 ? _989 : _988;
    assign _979 = ~ PHASE_11;
    assign read_enable_42 = _102 & _979;
    assign data_49 = wr_d3;
    assign _976 = _137[5:5];
    assign _975 = _137[4:4];
    assign _974 = _137[3:3];
    assign _973 = _137[2:2];
    assign _972 = _137[1:1];
    assign _971 = _137[0:0];
    assign _977 = { _971, _972, _973, _974, _975, _976 };
    assign address_53 = PHASE_11 ? _60 : _977;
    assign _968 = ~ PHASE_11;
    assign read_enable_43 = _102 & _968;
    assign _966 = _62[3:3];
    assign write_enable_53 = _966 & PHASE_11;
    assign _970 = write_enable_53 | read_enable_43;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_25
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_970), .regcea(vdd), .wea(write_enable_53), .addra(address_53), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_42), .regceb(vdd), .web(write_enable_52), .addrb(address_52), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_993[131:131]), .sbiterrb(_993[130:130]), .doutb(_993[129:66]), .dbiterra(_993[65:65]), .sbiterra(_993[64:64]), .douta(_993[63:0]) );
    assign _994 = _993[63:0];
    assign _927 = ~ PHASE_11;
    assign _35 = _927;
    always @(posedge _84) begin
        if (_82)
            PHASE_11 <= _925;
        else
            if (_72)
                PHASE_11 <= _35;
    end
    assign _1008 = PHASE_11 ? _1007 : _994;
    assign address_54 = _951 ? _199 : _172;
    assign _958 = ~ _951;
    assign read_enable_44 = _102 & _958;
    assign write_enable_54 = _942 & _951;
    assign _960 = write_enable_54 | read_enable_44;
    assign address_55 = _951 ? _164 : _137;
    assign _953 = ~ _951;
    assign read_enable_45 = _102 & _953;
    assign _951 = ~ PHASE_12;
    assign write_enable_55 = _935 & _951;
    assign _955 = write_enable_55 | read_enable_45;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_26
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_955), .regcea(vdd), .wea(write_enable_55), .addra(address_55), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_960), .regceb(vdd), .web(write_enable_54), .addrb(address_54), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_963[131:131]), .sbiterrb(_963[130:130]), .doutb(_963[129:66]), .dbiterra(_963[65:65]), .sbiterra(_963[64:64]), .douta(_963[63:0]) );
    assign _964 = _963[63:0];
    assign _1019 = _1018[127:64];
    assign data_51 = _1019;
    assign address_56 = PHASE_12 ? _199 : _172;
    assign _944 = ~ PHASE_12;
    assign read_enable_46 = _102 & _944;
    assign _941 = ~ _130;
    assign _942 = _129 & _941;
    assign write_enable_56 = _942 & PHASE_12;
    assign _946 = write_enable_56 | read_enable_46;
    assign address_57 = PHASE_12 ? _164 : _137;
    assign _937 = ~ PHASE_12;
    assign read_enable_47 = _102 & _937;
    assign _934 = ~ _130;
    assign _935 = _129 & _934;
    assign write_enable_57 = _935 & PHASE_12;
    assign _939 = write_enable_57 | read_enable_47;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_27
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_939), .regcea(vdd), .wea(write_enable_57), .addra(address_57), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_946), .regceb(vdd), .web(write_enable_56), .addrb(address_56), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_949[131:131]), .sbiterrb(_949[130:130]), .doutb(_949[129:66]), .dbiterra(_949[65:65]), .sbiterra(_949[64:64]), .douta(_949[63:0]) );
    assign _950 = _949[63:0];
    assign _1020 = ~ PHASE_12;
    assign _37 = _1020;
    always @(posedge _84) begin
        if (_82)
            PHASE_12 <= _932;
        else
            if (_99)
                PHASE_12 <= _37;
    end
    assign q0_3 = PHASE_12 ? _964 : _950;
    always @(posedge _84) begin
        if (_82)
            _930 <= _929;
        else
            _930 <= _92;
    end
    assign _1009 = _930 ? _1008 : q0_3;
    dp_26
        dp_2
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1009), .d2(_1016), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_1018[191:128]), .q2(_1018[127:64]), .q1(_1018[63:0]) );
    assign _1021 = _1018[63:0];
    assign data_55 = _1021;
    assign address_58 = PHASE_13 ? _164 : _68;
    assign _1085 = ~ PHASE_13;
    assign _1084 = _70[3:3];
    assign read_enable_48 = _1084 & _1085;
    always @(posedge _84) begin
        if (_82)
            _1055 <= _1054;
        else
            _1055 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _1058 <= _1057;
        else
            _1058 <= _1055;
    end
    always @(posedge _84) begin
        if (_82)
            _1061 <= _1060;
        else
            _1061 <= _1058;
    end
    always @(posedge _84) begin
        if (_82)
            _1064 <= _1063;
        else
            _1064 <= _1061;
    end
    always @(posedge _84) begin
        if (_82)
            _1067 <= _1066;
        else
            _1067 <= _1064;
    end
    always @(posedge _84) begin
        if (_82)
            _1070 <= _1069;
        else
            _1070 <= _1067;
    end
    always @(posedge _84) begin
        if (_82)
            _1073 <= _1072;
        else
            _1073 <= _1070;
    end
    always @(posedge _84) begin
        if (_82)
            _1076 <= _1075;
        else
            _1076 <= _1073;
    end
    always @(posedge _84) begin
        if (_82)
            _1079 <= _1078;
        else
            _1079 <= _1076;
    end
    assign _1080 = ~ _1079;
    always @(posedge _84) begin
        if (_82)
            _1028 <= _1027;
        else
            _1028 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1031 <= _1030;
        else
            _1031 <= _1028;
    end
    always @(posedge _84) begin
        if (_82)
            _1034 <= _1033;
        else
            _1034 <= _1031;
    end
    always @(posedge _84) begin
        if (_82)
            _1037 <= _1036;
        else
            _1037 <= _1034;
    end
    always @(posedge _84) begin
        if (_82)
            _1040 <= _1039;
        else
            _1040 <= _1037;
    end
    always @(posedge _84) begin
        if (_82)
            _1043 <= _1042;
        else
            _1043 <= _1040;
    end
    always @(posedge _84) begin
        if (_82)
            _1046 <= _1045;
        else
            _1046 <= _1043;
    end
    always @(posedge _84) begin
        if (_82)
            _1049 <= _1048;
        else
            _1049 <= _1046;
    end
    always @(posedge _84) begin
        if (_82)
            _1052 <= _1051;
        else
            _1052 <= _1049;
    end
    assign _1081 = _1052 & _1080;
    assign _1082 = _129 & _1081;
    assign write_enable_58 = _1082 & PHASE_13;
    assign _1087 = write_enable_58 | read_enable_48;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_28
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1087), .regcea(vdd), .wea(write_enable_58), .addra(address_58), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_49), .regceb(vdd), .web(write_enable_49), .addrb(address_49), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1094[131:131]), .sbiterrb(_1094[130:130]), .doutb(_1094[129:66]), .dbiterra(_1094[65:65]), .sbiterra(_1094[64:64]), .douta(_1094[63:0]) );
    assign _1095 = _1094[63:0];
    assign _1025 = ~ PHASE_13;
    assign _39 = _1025;
    always @(posedge _84) begin
        if (_82)
            PHASE_13 <= _1023;
        else
            if (_72)
                PHASE_13 <= _39;
    end
    assign _1107 = PHASE_13 ? _1106 : _1095;
    assign address_59 = _1280 ? _199 : _1275;
    assign write_enable_59 = _1273 & _1280;
    assign address_60 = _1280 ? _164 : _68;
    assign _1282 = ~ _1280;
    assign read_enable_49 = _1268 & _1282;
    assign _1280 = ~ PHASE_16;
    assign write_enable_60 = _1266 & _1280;
    assign _1284 = write_enable_60 | read_enable_49;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_29
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1284), .regcea(vdd), .wea(write_enable_60), .addra(address_60), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_59), .regceb(vdd), .web(write_enable_59), .addrb(address_59), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1289[131:131]), .sbiterrb(_1289[130:130]), .doutb(_1289[129:66]), .dbiterra(_1289[65:65]), .sbiterra(_1289[64:64]), .douta(_1289[63:0]) );
    assign _1290 = _1289[63:0];
    assign address_61 = PHASE_16 ? _199 : _1275;
    assign _1273 = _129 & _1236;
    assign write_enable_61 = _1273 & PHASE_16;
    assign _1198 = _1190[129:66];
    assign _1197 = _1177[129:66];
    assign _1199 = PHASE_14 ? _1198 : _1197;
    assign _1195 = _1147[129:66];
    assign _1194 = _1133[129:66];
    assign q1_4 = PHASE_15 ? _1195 : _1194;
    assign _1200 = _1114 ? _1199 : q1_4;
    assign address_62 = _1179 ? _1173 : _1172;
    assign _1185 = ~ _1179;
    assign read_enable_50 = _102 & _1185;
    assign address_63 = _1179 ? _60 : _1161;
    assign _1181 = ~ _1179;
    assign read_enable_51 = _102 & _1181;
    assign _1179 = ~ PHASE_14;
    assign write_enable_63 = _1150 & _1179;
    assign _1183 = write_enable_63 | read_enable_51;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_30
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1183), .regcea(vdd), .wea(write_enable_63), .addra(address_63), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_50), .regceb(vdd), .web(write_enable_62), .addrb(address_62), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1190[131:131]), .sbiterrb(_1190[130:130]), .doutb(_1190[129:66]), .dbiterra(_1190[65:65]), .sbiterra(_1190[64:64]), .douta(_1190[63:0]) );
    assign _1191 = _1190[63:0];
    assign _1171 = _172[5:5];
    assign _1170 = _172[4:4];
    assign _1169 = _172[3:3];
    assign _1168 = _172[2:2];
    assign _1167 = _172[1:1];
    assign _1166 = _172[0:0];
    assign _1172 = { _1166, _1167, _1168, _1169, _1170, _1171 };
    assign address_64 = PHASE_14 ? _1173 : _1172;
    assign _1163 = ~ PHASE_14;
    assign read_enable_52 = _102 & _1163;
    assign data_61 = wr_d2;
    assign _1160 = _137[5:5];
    assign _1159 = _137[4:4];
    assign _1158 = _137[3:3];
    assign _1157 = _137[2:2];
    assign _1156 = _137[1:1];
    assign _1155 = _137[0:0];
    assign _1161 = { _1155, _1156, _1157, _1158, _1159, _1160 };
    assign address_65 = PHASE_14 ? _60 : _1161;
    assign _1152 = ~ PHASE_14;
    assign read_enable_53 = _102 & _1152;
    assign _1150 = _62[2:2];
    assign write_enable_65 = _1150 & PHASE_14;
    assign _1154 = write_enable_65 | read_enable_53;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_31
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1154), .regcea(vdd), .wea(write_enable_65), .addra(address_65), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_52), .regceb(vdd), .web(write_enable_64), .addrb(address_64), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1177[131:131]), .sbiterrb(_1177[130:130]), .doutb(_1177[129:66]), .dbiterra(_1177[65:65]), .sbiterra(_1177[64:64]), .douta(_1177[63:0]) );
    assign _1178 = _1177[63:0];
    assign _1111 = ~ PHASE_14;
    assign _43 = _1111;
    always @(posedge _84) begin
        if (_82)
            PHASE_14 <= _1109;
        else
            if (_72)
                PHASE_14 <= _43;
    end
    assign _1192 = PHASE_14 ? _1191 : _1178;
    assign address_66 = _1135 ? _199 : _172;
    assign _1142 = ~ _1135;
    assign read_enable_54 = _102 & _1142;
    assign write_enable_66 = _1126 & _1135;
    assign _1144 = write_enable_66 | read_enable_54;
    assign address_67 = _1135 ? _164 : _137;
    assign _1137 = ~ _1135;
    assign read_enable_55 = _102 & _1137;
    assign _1135 = ~ PHASE_15;
    assign write_enable_67 = _1119 & _1135;
    assign _1139 = write_enable_67 | read_enable_55;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_32
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1139), .regcea(vdd), .wea(write_enable_67), .addra(address_67), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1144), .regceb(vdd), .web(write_enable_66), .addrb(address_66), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1147[131:131]), .sbiterrb(_1147[130:130]), .doutb(_1147[129:66]), .dbiterra(_1147[65:65]), .sbiterra(_1147[64:64]), .douta(_1147[63:0]) );
    assign _1148 = _1147[63:0];
    assign _1203 = _1202[127:64];
    assign data_63 = _1203;
    assign address_68 = PHASE_15 ? _199 : _172;
    assign _1128 = ~ PHASE_15;
    assign read_enable_56 = _102 & _1128;
    assign _1125 = ~ _130;
    assign _1126 = _129 & _1125;
    assign write_enable_68 = _1126 & PHASE_15;
    assign _1130 = write_enable_68 | read_enable_56;
    assign address_69 = PHASE_15 ? _164 : _137;
    assign _1121 = ~ PHASE_15;
    assign read_enable_57 = _102 & _1121;
    assign _1118 = ~ _130;
    assign _1119 = _129 & _1118;
    assign write_enable_69 = _1119 & PHASE_15;
    assign _1123 = write_enable_69 | read_enable_57;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_33
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1123), .regcea(vdd), .wea(write_enable_69), .addra(address_69), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1130), .regceb(vdd), .web(write_enable_68), .addrb(address_68), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1133[131:131]), .sbiterrb(_1133[130:130]), .doutb(_1133[129:66]), .dbiterra(_1133[65:65]), .sbiterra(_1133[64:64]), .douta(_1133[63:0]) );
    assign _1134 = _1133[63:0];
    assign _1204 = ~ PHASE_15;
    assign _45 = _1204;
    always @(posedge _84) begin
        if (_82)
            PHASE_15 <= _1116;
        else
            if (_99)
                PHASE_15 <= _45;
    end
    assign q0_4 = PHASE_15 ? _1148 : _1134;
    always @(posedge _84) begin
        if (_82)
            _1114 <= _1113;
        else
            _1114 <= _92;
    end
    assign _1193 = _1114 ? _1192 : q0_4;
    dp_25
        dp_1
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1193), .d2(_1200), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_1202[191:128]), .q2(_1202[127:64]), .q1(_1202[63:0]) );
    assign _1205 = _1202[63:0];
    assign data_67 = _1205;
    assign address_70 = PHASE_16 ? _164 : _68;
    assign _1269 = ~ PHASE_16;
    assign _1268 = _70[2:2];
    assign read_enable_58 = _1268 & _1269;
    always @(posedge _84) begin
        if (_82)
            _1239 <= _1238;
        else
            _1239 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _1242 <= _1241;
        else
            _1242 <= _1239;
    end
    always @(posedge _84) begin
        if (_82)
            _1245 <= _1244;
        else
            _1245 <= _1242;
    end
    always @(posedge _84) begin
        if (_82)
            _1248 <= _1247;
        else
            _1248 <= _1245;
    end
    always @(posedge _84) begin
        if (_82)
            _1251 <= _1250;
        else
            _1251 <= _1248;
    end
    always @(posedge _84) begin
        if (_82)
            _1254 <= _1253;
        else
            _1254 <= _1251;
    end
    always @(posedge _84) begin
        if (_82)
            _1257 <= _1256;
        else
            _1257 <= _1254;
    end
    always @(posedge _84) begin
        if (_82)
            _1260 <= _1259;
        else
            _1260 <= _1257;
    end
    always @(posedge _84) begin
        if (_82)
            _1263 <= _1262;
        else
            _1263 <= _1260;
    end
    assign _1264 = ~ _1263;
    always @(posedge _84) begin
        if (_82)
            _1212 <= _1211;
        else
            _1212 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1215 <= _1214;
        else
            _1215 <= _1212;
    end
    always @(posedge _84) begin
        if (_82)
            _1218 <= _1217;
        else
            _1218 <= _1215;
    end
    always @(posedge _84) begin
        if (_82)
            _1221 <= _1220;
        else
            _1221 <= _1218;
    end
    always @(posedge _84) begin
        if (_82)
            _1224 <= _1223;
        else
            _1224 <= _1221;
    end
    always @(posedge _84) begin
        if (_82)
            _1227 <= _1226;
        else
            _1227 <= _1224;
    end
    always @(posedge _84) begin
        if (_82)
            _1230 <= _1229;
        else
            _1230 <= _1227;
    end
    always @(posedge _84) begin
        if (_82)
            _1233 <= _1232;
        else
            _1233 <= _1230;
    end
    always @(posedge _84) begin
        if (_82)
            _1236 <= _1235;
        else
            _1236 <= _1233;
    end
    assign _1265 = _1236 & _1264;
    assign _1266 = _129 & _1265;
    assign write_enable_70 = _1266 & PHASE_16;
    assign _1271 = write_enable_70 | read_enable_58;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_34
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1271), .regcea(vdd), .wea(write_enable_70), .addra(address_70), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_61), .regceb(vdd), .web(write_enable_61), .addrb(address_61), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1278[131:131]), .sbiterrb(_1278[130:130]), .doutb(_1278[129:66]), .dbiterra(_1278[65:65]), .sbiterra(_1278[64:64]), .douta(_1278[63:0]) );
    assign _1279 = _1278[63:0];
    assign _1209 = ~ PHASE_16;
    assign _47 = _1209;
    always @(posedge _84) begin
        if (_82)
            PHASE_16 <= _1207;
        else
            if (_72)
                PHASE_16 <= _47;
    end
    assign _1291 = PHASE_16 ? _1290 : _1279;
    assign address_71 = _1464 ? _199 : _1459;
    assign write_enable_71 = _1457 & _1464;
    assign address_72 = _1464 ? _164 : _68;
    assign _1466 = ~ _1464;
    assign read_enable_59 = _1452 & _1466;
    assign _1464 = ~ PHASE_19;
    assign write_enable_72 = _1450 & _1464;
    assign _1468 = write_enable_72 | read_enable_59;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_35
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1468), .regcea(vdd), .wea(write_enable_72), .addra(address_72), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_71), .regceb(vdd), .web(write_enable_71), .addrb(address_71), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1473[131:131]), .sbiterrb(_1473[130:130]), .doutb(_1473[129:66]), .dbiterra(_1473[65:65]), .sbiterra(_1473[64:64]), .douta(_1473[63:0]) );
    assign _1474 = _1473[63:0];
    assign address_73 = PHASE_19 ? _199 : _1459;
    assign _1457 = _129 & _1420;
    assign write_enable_73 = _1457 & PHASE_19;
    assign _1382 = _1374[129:66];
    assign _1381 = _1361[129:66];
    assign _1383 = PHASE_17 ? _1382 : _1381;
    assign _1379 = _1331[129:66];
    assign _1378 = _1317[129:66];
    assign q1_5 = PHASE_18 ? _1379 : _1378;
    assign _1384 = _1298 ? _1383 : q1_5;
    assign address_74 = _1363 ? _1357 : _1356;
    assign _1369 = ~ _1363;
    assign read_enable_60 = _102 & _1369;
    assign address_75 = _1363 ? _60 : _1345;
    assign _1365 = ~ _1363;
    assign read_enable_61 = _102 & _1365;
    assign _1363 = ~ PHASE_17;
    assign write_enable_75 = _1334 & _1363;
    assign _1367 = write_enable_75 | read_enable_61;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_36
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1367), .regcea(vdd), .wea(write_enable_75), .addra(address_75), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_60), .regceb(vdd), .web(write_enable_74), .addrb(address_74), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1374[131:131]), .sbiterrb(_1374[130:130]), .doutb(_1374[129:66]), .dbiterra(_1374[65:65]), .sbiterra(_1374[64:64]), .douta(_1374[63:0]) );
    assign _1375 = _1374[63:0];
    assign _1355 = _172[5:5];
    assign _1354 = _172[4:4];
    assign _1353 = _172[3:3];
    assign _1352 = _172[2:2];
    assign _1351 = _172[1:1];
    assign _1350 = _172[0:0];
    assign _1356 = { _1350, _1351, _1352, _1353, _1354, _1355 };
    assign address_76 = PHASE_17 ? _1357 : _1356;
    assign _1347 = ~ PHASE_17;
    assign read_enable_62 = _102 & _1347;
    assign data_73 = wr_d1;
    assign _1344 = _137[5:5];
    assign _1343 = _137[4:4];
    assign _1342 = _137[3:3];
    assign _1341 = _137[2:2];
    assign _1340 = _137[1:1];
    assign _1339 = _137[0:0];
    assign _1345 = { _1339, _1340, _1341, _1342, _1343, _1344 };
    assign address_77 = PHASE_17 ? _60 : _1345;
    assign _1336 = ~ PHASE_17;
    assign read_enable_63 = _102 & _1336;
    assign _1334 = _62[1:1];
    assign write_enable_77 = _1334 & PHASE_17;
    assign _1338 = write_enable_77 | read_enable_63;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_37
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1338), .regcea(vdd), .wea(write_enable_77), .addra(address_77), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_62), .regceb(vdd), .web(write_enable_76), .addrb(address_76), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1361[131:131]), .sbiterrb(_1361[130:130]), .doutb(_1361[129:66]), .dbiterra(_1361[65:65]), .sbiterra(_1361[64:64]), .douta(_1361[63:0]) );
    assign _1362 = _1361[63:0];
    assign _1295 = ~ PHASE_17;
    assign _51 = _1295;
    always @(posedge _84) begin
        if (_82)
            PHASE_17 <= _1293;
        else
            if (_72)
                PHASE_17 <= _51;
    end
    assign _1376 = PHASE_17 ? _1375 : _1362;
    assign address_78 = _1319 ? _199 : _172;
    assign _1326 = ~ _1319;
    assign read_enable_64 = _102 & _1326;
    assign write_enable_78 = _1310 & _1319;
    assign _1328 = write_enable_78 | read_enable_64;
    assign address_79 = _1319 ? _164 : _137;
    assign _1321 = ~ _1319;
    assign read_enable_65 = _102 & _1321;
    assign _1319 = ~ PHASE_18;
    assign write_enable_79 = _1303 & _1319;
    assign _1323 = write_enable_79 | read_enable_65;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_38
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1323), .regcea(vdd), .wea(write_enable_79), .addra(address_79), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1328), .regceb(vdd), .web(write_enable_78), .addrb(address_78), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1331[131:131]), .sbiterrb(_1331[130:130]), .doutb(_1331[129:66]), .dbiterra(_1331[65:65]), .sbiterra(_1331[64:64]), .douta(_1331[63:0]) );
    assign _1332 = _1331[63:0];
    assign _1387 = _1386[127:64];
    assign data_75 = _1387;
    assign address_80 = PHASE_18 ? _199 : _172;
    assign _1312 = ~ PHASE_18;
    assign read_enable_66 = _102 & _1312;
    assign _1309 = ~ _130;
    assign _1310 = _129 & _1309;
    assign write_enable_80 = _1310 & PHASE_18;
    assign _1314 = write_enable_80 | read_enable_66;
    assign address_81 = PHASE_18 ? _164 : _137;
    assign _1305 = ~ PHASE_18;
    assign read_enable_67 = _102 & _1305;
    assign _1302 = ~ _130;
    assign _1303 = _129 & _1302;
    assign write_enable_81 = _1303 & PHASE_18;
    assign _1307 = write_enable_81 | read_enable_67;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_39
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1307), .regcea(vdd), .wea(write_enable_81), .addra(address_81), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1314), .regceb(vdd), .web(write_enable_80), .addrb(address_80), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1317[131:131]), .sbiterrb(_1317[130:130]), .doutb(_1317[129:66]), .dbiterra(_1317[65:65]), .sbiterra(_1317[64:64]), .douta(_1317[63:0]) );
    assign _1318 = _1317[63:0];
    assign _1388 = ~ PHASE_18;
    assign _53 = _1388;
    always @(posedge _84) begin
        if (_82)
            PHASE_18 <= _1300;
        else
            if (_99)
                PHASE_18 <= _53;
    end
    assign q0_5 = PHASE_18 ? _1332 : _1318;
    always @(posedge _84) begin
        if (_82)
            _1298 <= _1297;
        else
            _1298 <= _92;
    end
    assign _1377 = _1298 ? _1376 : q0_5;
    dp_24
        dp_0
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1377), .d2(_1384), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_1386[191:128]), .q2(_1386[127:64]), .q1(_1386[63:0]) );
    assign _1389 = _1386[63:0];
    assign data_79 = _1389;
    assign address_82 = PHASE_19 ? _164 : _68;
    assign _1453 = ~ PHASE_19;
    assign _1452 = _70[1:1];
    assign read_enable_68 = _1452 & _1453;
    always @(posedge _84) begin
        if (_82)
            _1423 <= _1422;
        else
            _1423 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _1426 <= _1425;
        else
            _1426 <= _1423;
    end
    always @(posedge _84) begin
        if (_82)
            _1429 <= _1428;
        else
            _1429 <= _1426;
    end
    always @(posedge _84) begin
        if (_82)
            _1432 <= _1431;
        else
            _1432 <= _1429;
    end
    always @(posedge _84) begin
        if (_82)
            _1435 <= _1434;
        else
            _1435 <= _1432;
    end
    always @(posedge _84) begin
        if (_82)
            _1438 <= _1437;
        else
            _1438 <= _1435;
    end
    always @(posedge _84) begin
        if (_82)
            _1441 <= _1440;
        else
            _1441 <= _1438;
    end
    always @(posedge _84) begin
        if (_82)
            _1444 <= _1443;
        else
            _1444 <= _1441;
    end
    always @(posedge _84) begin
        if (_82)
            _1447 <= _1446;
        else
            _1447 <= _1444;
    end
    assign _1448 = ~ _1447;
    always @(posedge _84) begin
        if (_82)
            _1396 <= _1395;
        else
            _1396 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1399 <= _1398;
        else
            _1399 <= _1396;
    end
    always @(posedge _84) begin
        if (_82)
            _1402 <= _1401;
        else
            _1402 <= _1399;
    end
    always @(posedge _84) begin
        if (_82)
            _1405 <= _1404;
        else
            _1405 <= _1402;
    end
    always @(posedge _84) begin
        if (_82)
            _1408 <= _1407;
        else
            _1408 <= _1405;
    end
    always @(posedge _84) begin
        if (_82)
            _1411 <= _1410;
        else
            _1411 <= _1408;
    end
    always @(posedge _84) begin
        if (_82)
            _1414 <= _1413;
        else
            _1414 <= _1411;
    end
    always @(posedge _84) begin
        if (_82)
            _1417 <= _1416;
        else
            _1417 <= _1414;
    end
    always @(posedge _84) begin
        if (_82)
            _1420 <= _1419;
        else
            _1420 <= _1417;
    end
    assign _1449 = _1420 & _1448;
    assign _1450 = _129 & _1449;
    assign write_enable_82 = _1450 & PHASE_19;
    assign _1455 = write_enable_82 | read_enable_68;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_40
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1455), .regcea(vdd), .wea(write_enable_82), .addra(address_82), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_73), .regceb(vdd), .web(write_enable_73), .addrb(address_73), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1462[131:131]), .sbiterrb(_1462[130:130]), .doutb(_1462[129:66]), .dbiterra(_1462[65:65]), .sbiterra(_1462[64:64]), .douta(_1462[63:0]) );
    assign _1463 = _1462[63:0];
    assign _1393 = ~ PHASE_19;
    assign _55 = _1393;
    always @(posedge _84) begin
        if (_82)
            PHASE_19 <= _1391;
        else
            if (_72)
                PHASE_19 <= _55;
    end
    assign _1475 = PHASE_19 ? _1474 : _1463;
    assign address_83 = _1648 ? _199 : _1643;
    assign write_enable_83 = _1641 & _1648;
    assign address_84 = _1648 ? _164 : _68;
    assign _1650 = ~ _1648;
    assign read_enable_69 = _1636 & _1650;
    assign _1648 = ~ PHASE_22;
    assign write_enable_84 = _1634 & _1648;
    assign _1652 = write_enable_84 | read_enable_69;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_41
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1652), .regcea(vdd), .wea(write_enable_84), .addra(address_84), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_83), .regceb(vdd), .web(write_enable_83), .addrb(address_83), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1657[131:131]), .sbiterrb(_1657[130:130]), .doutb(_1657[129:66]), .dbiterra(_1657[65:65]), .sbiterra(_1657[64:64]), .douta(_1657[63:0]) );
    assign _1658 = _1657[63:0];
    assign address_85 = PHASE_22 ? _199 : _1643;
    assign _1641 = _129 & _1604;
    assign write_enable_85 = _1641 & PHASE_22;
    assign _280 = _91[490:487];
    assign _279 = _91[486:486];
    assign _277 = _91[482:482];
    assign _276 = _91[481:418];
    assign _275 = _91[417:354];
    assign _274 = _91[353:290];
    assign _273 = _91[289:226];
    assign _272 = _91[225:162];
    assign _271 = _91[161:98];
    assign _270 = _91[97:34];
    assign _1566 = _1558[129:66];
    assign _1565 = _1545[129:66];
    assign _1567 = PHASE_20 ? _1566 : _1565;
    assign _1563 = _1515[129:66];
    assign _1562 = _1501[129:66];
    assign q1_6 = PHASE_21 ? _1563 : _1562;
    assign _1568 = _1482 ? _1567 : q1_6;
    assign address_86 = _1547 ? _1541 : _1540;
    assign _1553 = ~ _1547;
    assign read_enable_70 = _102 & _1553;
    assign address_87 = _1547 ? _60 : _1529;
    assign _1549 = ~ _1547;
    assign read_enable_71 = _102 & _1549;
    assign _1547 = ~ PHASE_20;
    assign write_enable_87 = _1518 & _1547;
    assign _1551 = write_enable_87 | read_enable_71;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_42
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1551), .regcea(vdd), .wea(write_enable_87), .addra(address_87), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_70), .regceb(vdd), .web(write_enable_86), .addrb(address_86), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1558[131:131]), .sbiterrb(_1558[130:130]), .doutb(_1558[129:66]), .dbiterra(_1558[65:65]), .sbiterra(_1558[64:64]), .douta(_1558[63:0]) );
    assign _1559 = _1558[63:0];
    assign _1539 = _172[5:5];
    assign _1538 = _172[4:4];
    assign _1537 = _172[3:3];
    assign _1536 = _172[2:2];
    assign _1535 = _172[1:1];
    assign _1534 = _172[0:0];
    assign _1540 = { _1534, _1535, _1536, _1537, _1538, _1539 };
    assign address_88 = PHASE_20 ? _1541 : _1540;
    assign _1531 = ~ PHASE_20;
    assign read_enable_72 = _102 & _1531;
    assign data_85 = wr_d0;
    assign _60 = wr_addr;
    assign _1528 = _137[5:5];
    assign _1527 = _137[4:4];
    assign _1526 = _137[3:3];
    assign _1525 = _137[2:2];
    assign _1524 = _137[1:1];
    assign _1523 = _137[0:0];
    assign _1529 = { _1523, _1524, _1525, _1526, _1527, _1528 };
    assign address_89 = PHASE_20 ? _60 : _1529;
    assign _1520 = ~ PHASE_20;
    assign read_enable_73 = _102 & _1520;
    assign _62 = wr_en;
    assign _1518 = _62[0:0];
    assign write_enable_89 = _1518 & PHASE_20;
    assign _1522 = write_enable_89 | read_enable_73;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_43
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1522), .regcea(vdd), .wea(write_enable_89), .addra(address_89), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_72), .regceb(vdd), .web(write_enable_88), .addrb(address_88), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1545[131:131]), .sbiterrb(_1545[130:130]), .doutb(_1545[129:66]), .dbiterra(_1545[65:65]), .sbiterra(_1545[64:64]), .douta(_1545[63:0]) );
    assign _1546 = _1545[63:0];
    assign _1479 = ~ PHASE_20;
    assign _63 = _1479;
    always @(posedge _84) begin
        if (_82)
            PHASE_20 <= _1477;
        else
            if (_72)
                PHASE_20 <= _63;
    end
    assign _1560 = PHASE_20 ? _1559 : _1546;
    assign address_90 = _1503 ? _199 : _172;
    assign _1510 = ~ _1503;
    assign read_enable_74 = _102 & _1510;
    assign write_enable_90 = _1494 & _1503;
    assign _1512 = write_enable_90 | read_enable_74;
    assign address_91 = _1503 ? _164 : _137;
    assign _1505 = ~ _1503;
    assign read_enable_75 = _102 & _1505;
    assign _1503 = ~ PHASE_21;
    assign write_enable_91 = _1487 & _1503;
    assign _1507 = write_enable_91 | read_enable_75;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_44
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1507), .regcea(vdd), .wea(write_enable_91), .addra(address_91), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1512), .regceb(vdd), .web(write_enable_90), .addrb(address_90), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1515[131:131]), .sbiterrb(_1515[130:130]), .doutb(_1515[129:66]), .dbiterra(_1515[65:65]), .sbiterra(_1515[64:64]), .douta(_1515[63:0]) );
    assign _1516 = _1515[63:0];
    assign _1571 = _1570[127:64];
    assign data_87 = _1571;
    always @(posedge _84) begin
        if (_82)
            _175 <= _174;
        else
            _175 <= _172;
    end
    always @(posedge _84) begin
        if (_82)
            _178 <= _177;
        else
            _178 <= _175;
    end
    always @(posedge _84) begin
        if (_82)
            _181 <= _180;
        else
            _181 <= _178;
    end
    always @(posedge _84) begin
        if (_82)
            _184 <= _183;
        else
            _184 <= _181;
    end
    always @(posedge _84) begin
        if (_82)
            _187 <= _186;
        else
            _187 <= _184;
    end
    always @(posedge _84) begin
        if (_82)
            _190 <= _189;
        else
            _190 <= _187;
    end
    always @(posedge _84) begin
        if (_82)
            _193 <= _192;
        else
            _193 <= _190;
    end
    always @(posedge _84) begin
        if (_82)
            _196 <= _195;
        else
            _196 <= _193;
    end
    always @(posedge _84) begin
        if (_82)
            _199 <= _198;
        else
            _199 <= _196;
    end
    assign _172 = _91[33:28];
    assign address_92 = PHASE_21 ? _199 : _172;
    assign _1496 = ~ PHASE_21;
    assign read_enable_76 = _102 & _1496;
    assign _1493 = ~ _130;
    assign _1494 = _129 & _1493;
    assign write_enable_92 = _1494 & PHASE_21;
    assign _1498 = write_enable_92 | read_enable_76;
    assign address_93 = PHASE_21 ? _164 : _137;
    assign _1489 = ~ PHASE_21;
    assign read_enable_77 = _102 & _1489;
    assign _1486 = ~ _130;
    assign _1487 = _129 & _1486;
    assign write_enable_93 = _1487 & PHASE_21;
    assign _1491 = write_enable_93 | read_enable_77;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_45
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1491), .regcea(vdd), .wea(write_enable_93), .addra(address_93), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1498), .regceb(vdd), .web(write_enable_92), .addrb(address_92), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1501[131:131]), .sbiterrb(_1501[130:130]), .doutb(_1501[129:66]), .dbiterra(_1501[65:65]), .sbiterra(_1501[64:64]), .douta(_1501[63:0]) );
    assign _1502 = _1501[63:0];
    assign _99 = _91[492:492];
    assign _1572 = ~ PHASE_21;
    assign _65 = _1572;
    always @(posedge _84) begin
        if (_82)
            PHASE_21 <= _1484;
        else
            if (_99)
                PHASE_21 <= _65;
    end
    assign q0_6 = PHASE_21 ? _1516 : _1502;
    assign _92 = _91[483:483];
    always @(posedge _84) begin
        if (_82)
            _1482 <= _1481;
        else
            _1482 <= _92;
    end
    assign _1561 = _1482 ? _1560 : q0_6;
    dp_23
        dp
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1561), .d2(_1568), .omegas0(_270), .omegas1(_271), .omegas2(_272), .omegas3(_273), .omegas4(_274), .omegas5(_275), .omegas6(_276), .start_twiddles(_277), .twiddle_stage(_278), .valid(_279), .index(_280), .twiddle_update_q(_1570[191:128]), .q2(_1570[127:64]), .q1(_1570[63:0]) );
    assign _1573 = _1570[63:0];
    assign data_91 = _1573;
    assign _137 = _91[27:22];
    always @(posedge _84) begin
        if (_82)
            _140 <= _139;
        else
            _140 <= _137;
    end
    always @(posedge _84) begin
        if (_82)
            _143 <= _142;
        else
            _143 <= _140;
    end
    always @(posedge _84) begin
        if (_82)
            _146 <= _145;
        else
            _146 <= _143;
    end
    always @(posedge _84) begin
        if (_82)
            _149 <= _148;
        else
            _149 <= _146;
    end
    always @(posedge _84) begin
        if (_82)
            _152 <= _151;
        else
            _152 <= _149;
    end
    always @(posedge _84) begin
        if (_82)
            _155 <= _154;
        else
            _155 <= _152;
    end
    always @(posedge _84) begin
        if (_82)
            _158 <= _157;
        else
            _158 <= _155;
    end
    always @(posedge _84) begin
        if (_82)
            _161 <= _160;
        else
            _161 <= _158;
    end
    always @(posedge _84) begin
        if (_82)
            _164 <= _163;
        else
            _164 <= _161;
    end
    assign _68 = rd_addr;
    assign address_94 = PHASE_22 ? _164 : _68;
    assign _1637 = ~ PHASE_22;
    assign _70 = rd_en;
    assign _1636 = _70[0:0];
    assign read_enable_78 = _1636 & _1637;
    assign _278 = _91[485:485];
    always @(posedge _84) begin
        if (_82)
            _1607 <= _1606;
        else
            _1607 <= _278;
    end
    always @(posedge _84) begin
        if (_82)
            _1610 <= _1609;
        else
            _1610 <= _1607;
    end
    always @(posedge _84) begin
        if (_82)
            _1613 <= _1612;
        else
            _1613 <= _1610;
    end
    always @(posedge _84) begin
        if (_82)
            _1616 <= _1615;
        else
            _1616 <= _1613;
    end
    always @(posedge _84) begin
        if (_82)
            _1619 <= _1618;
        else
            _1619 <= _1616;
    end
    always @(posedge _84) begin
        if (_82)
            _1622 <= _1621;
        else
            _1622 <= _1619;
    end
    always @(posedge _84) begin
        if (_82)
            _1625 <= _1624;
        else
            _1625 <= _1622;
    end
    always @(posedge _84) begin
        if (_82)
            _1628 <= _1627;
        else
            _1628 <= _1625;
    end
    always @(posedge _84) begin
        if (_82)
            _1631 <= _1630;
        else
            _1631 <= _1628;
    end
    assign _1632 = ~ _1631;
    assign _130 = _91[484:484];
    always @(posedge _84) begin
        if (_82)
            _1580 <= _1579;
        else
            _1580 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1583 <= _1582;
        else
            _1583 <= _1580;
    end
    always @(posedge _84) begin
        if (_82)
            _1586 <= _1585;
        else
            _1586 <= _1583;
    end
    always @(posedge _84) begin
        if (_82)
            _1589 <= _1588;
        else
            _1589 <= _1586;
    end
    always @(posedge _84) begin
        if (_82)
            _1592 <= _1591;
        else
            _1592 <= _1589;
    end
    always @(posedge _84) begin
        if (_82)
            _1595 <= _1594;
        else
            _1595 <= _1592;
    end
    always @(posedge _84) begin
        if (_82)
            _1598 <= _1597;
        else
            _1598 <= _1595;
    end
    always @(posedge _84) begin
        if (_82)
            _1601 <= _1600;
        else
            _1601 <= _1598;
    end
    always @(posedge _84) begin
        if (_82)
            _1604 <= _1603;
        else
            _1604 <= _1601;
    end
    assign _1633 = _1604 & _1632;
    assign _102 = _91[491:491];
    always @(posedge _84) begin
        if (_82)
            _105 <= _104;
        else
            _105 <= _102;
    end
    always @(posedge _84) begin
        if (_82)
            _108 <= _107;
        else
            _108 <= _105;
    end
    always @(posedge _84) begin
        if (_82)
            _111 <= _110;
        else
            _111 <= _108;
    end
    always @(posedge _84) begin
        if (_82)
            _114 <= _113;
        else
            _114 <= _111;
    end
    always @(posedge _84) begin
        if (_82)
            _117 <= _116;
        else
            _117 <= _114;
    end
    always @(posedge _84) begin
        if (_82)
            _120 <= _119;
        else
            _120 <= _117;
    end
    always @(posedge _84) begin
        if (_82)
            _123 <= _122;
        else
            _123 <= _120;
    end
    always @(posedge _84) begin
        if (_82)
            _126 <= _125;
        else
            _126 <= _123;
    end
    always @(posedge _84) begin
        if (_82)
            _129 <= _128;
        else
            _129 <= _126;
    end
    assign _1634 = _129 & _1633;
    assign write_enable_94 = _1634 & PHASE_22;
    assign _1639 = write_enable_94 | read_enable_78;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(4096), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(6), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(6), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_46
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1639), .regcea(vdd), .wea(write_enable_94), .addra(address_94), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_85), .regceb(vdd), .web(write_enable_85), .addrb(address_85), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1646[131:131]), .sbiterrb(_1646[130:130]), .doutb(_1646[129:66]), .dbiterra(_1646[65:65]), .sbiterra(_1646[64:64]), .douta(_1646[63:0]) );
    assign _1647 = _1646[63:0];
    assign _72 = flip;
    assign _1577 = ~ PHASE_22;
    assign _73 = _1577;
    always @(posedge _84) begin
        if (_82)
            PHASE_22 <= _1575;
        else
            if (_72)
                PHASE_22 <= _73;
    end
    assign _1659 = PHASE_22 ? _1658 : _1647;
    assign _76 = first_4step_pass;
    assign _78 = first_iter;
    assign _80 = start;
    assign _82 = clear;
    assign _84 = clock;
    ctrl
        ctrl
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .first_4step_pass(_76), .flip(_91[492:492]), .read_write_enable(_91[491:491]), .index(_91[490:487]), .valid(_91[486:486]), .twiddle_stage(_91[485:485]), .last_stage(_91[484:484]), .first_stage(_91[483:483]), .start_twiddles(_91[482:482]), .omegas6(_91[481:418]), .omegas5(_91[417:354]), .omegas4(_91[353:290]), .omegas3(_91[289:226]), .omegas2(_91[225:162]), .omegas1(_91[161:98]), .omegas0(_91[97:34]), .addr2(_91[33:28]), .addr1(_91[27:22]), .m(_91[21:16]), .k(_91[15:10]), .j(_91[9:4]), .i(_91[3:1]), .done_(_91[0:0]) );
    assign _1660 = _91[0:0];

    /* aliases */
    assign data_0 = data;
    assign data_2 = data_1;
    assign data_4 = data_3;
    assign data_5 = data_3;
    assign data_6 = data_3;
    assign data_8 = data_7;
    assign data_9 = data_7;
    assign data_10 = data_7;
    assign data_12 = data_11;
    assign data_14 = data_13;
    assign data_16 = data_15;
    assign data_17 = data_15;
    assign data_18 = data_15;
    assign data_20 = data_19;
    assign data_21 = data_19;
    assign data_22 = data_19;
    assign data_24 = data_23;
    assign data_26 = data_25;
    assign data_28 = data_27;
    assign data_29 = data_27;
    assign data_30 = data_27;
    assign data_32 = data_31;
    assign data_33 = data_31;
    assign data_34 = data_31;
    assign data_36 = data_35;
    assign data_38 = data_37;
    assign data_40 = data_39;
    assign data_41 = data_39;
    assign data_42 = data_39;
    assign data_44 = data_43;
    assign data_45 = data_43;
    assign data_46 = data_43;
    assign data_48 = data_47;
    assign data_50 = data_49;
    assign data_52 = data_51;
    assign data_53 = data_51;
    assign data_54 = data_51;
    assign data_56 = data_55;
    assign data_57 = data_55;
    assign data_58 = data_55;
    assign data_60 = data_59;
    assign data_62 = data_61;
    assign data_64 = data_63;
    assign data_65 = data_63;
    assign data_66 = data_63;
    assign data_68 = data_67;
    assign data_69 = data_67;
    assign data_70 = data_67;
    assign data_72 = data_71;
    assign data_74 = data_73;
    assign data_76 = data_75;
    assign data_77 = data_75;
    assign data_78 = data_75;
    assign data_80 = data_79;
    assign data_81 = data_79;
    assign data_82 = data_79;
    assign data_84 = data_83;
    assign data_86 = data_85;
    assign data_88 = data_87;
    assign data_89 = data_87;
    assign data_90 = data_87;
    assign data_92 = data_91;
    assign data_93 = data_91;
    assign data_94 = data_91;

    /* output assignments */
    assign done_ = _1660;
    assign rd_q0 = _1659;
    assign rd_q1 = _1475;
    assign rd_q2 = _1291;
    assign rd_q3 = _1107;
    assign rd_q4 = _923;
    assign rd_q5 = _739;
    assign rd_q6 = _555;
    assign rd_q7 = _371;

endmodule
module multi_parallel_cores (
    rd_addr3,
    wr_addr3,
    wr_d_3_7,
    wr_d_3_6,
    wr_d_3_5,
    wr_d_3_4,
    wr_d_3_3,
    wr_d_3_2,
    wr_d_3_1,
    wr_d_3_0,
    rd_addr2,
    wr_addr2,
    wr_d_2_7,
    wr_d_2_6,
    wr_d_2_5,
    wr_d_2_4,
    wr_d_2_3,
    wr_d_2_2,
    wr_d_2_1,
    wr_d_2_0,
    rd_addr1,
    wr_addr1,
    wr_d_1_7,
    wr_d_1_6,
    wr_d_1_5,
    wr_d_1_4,
    wr_d_1_3,
    wr_d_1_2,
    wr_d_1_1,
    wr_d_1_0,
    rd_addr0,
    rd_en,
    wr_addr0,
    wr_en,
    wr_d_0_7,
    wr_d_0_6,
    wr_d_0_5,
    wr_d_0_4,
    wr_d_0_3,
    wr_d_0_2,
    wr_d_0_1,
    wr_d_0_0,
    flip,
    first_iter,
    first_4step_pass,
    start,
    clear,
    clock,
    done_,
    rd_d_0_0,
    rd_d_0_1,
    rd_d_0_2,
    rd_d_0_3,
    rd_d_0_4,
    rd_d_0_5,
    rd_d_0_6,
    rd_d_0_7,
    rd_d_1_0,
    rd_d_1_1,
    rd_d_1_2,
    rd_d_1_3,
    rd_d_1_4,
    rd_d_1_5,
    rd_d_1_6,
    rd_d_1_7,
    rd_d_2_0,
    rd_d_2_1,
    rd_d_2_2,
    rd_d_2_3,
    rd_d_2_4,
    rd_d_2_5,
    rd_d_2_6,
    rd_d_2_7,
    rd_d_3_0,
    rd_d_3_1,
    rd_d_3_2,
    rd_d_3_3,
    rd_d_3_4,
    rd_d_3_5,
    rd_d_3_6,
    rd_d_3_7
);

    input [5:0] rd_addr3;
    input [5:0] wr_addr3;
    input [63:0] wr_d_3_7;
    input [63:0] wr_d_3_6;
    input [63:0] wr_d_3_5;
    input [63:0] wr_d_3_4;
    input [63:0] wr_d_3_3;
    input [63:0] wr_d_3_2;
    input [63:0] wr_d_3_1;
    input [63:0] wr_d_3_0;
    input [5:0] rd_addr2;
    input [5:0] wr_addr2;
    input [63:0] wr_d_2_7;
    input [63:0] wr_d_2_6;
    input [63:0] wr_d_2_5;
    input [63:0] wr_d_2_4;
    input [63:0] wr_d_2_3;
    input [63:0] wr_d_2_2;
    input [63:0] wr_d_2_1;
    input [63:0] wr_d_2_0;
    input [5:0] rd_addr1;
    input [5:0] wr_addr1;
    input [63:0] wr_d_1_7;
    input [63:0] wr_d_1_6;
    input [63:0] wr_d_1_5;
    input [63:0] wr_d_1_4;
    input [63:0] wr_d_1_3;
    input [63:0] wr_d_1_2;
    input [63:0] wr_d_1_1;
    input [63:0] wr_d_1_0;
    input [5:0] rd_addr0;
    input [3:0] rd_en;
    input [5:0] wr_addr0;
    input [3:0] wr_en;
    input [63:0] wr_d_0_7;
    input [63:0] wr_d_0_6;
    input [63:0] wr_d_0_5;
    input [63:0] wr_d_0_4;
    input [63:0] wr_d_0_3;
    input [63:0] wr_d_0_2;
    input [63:0] wr_d_0_1;
    input [63:0] wr_d_0_0;
    input flip;
    input first_iter;
    input first_4step_pass;
    input start;
    input clear;
    input clock;
    output done_;
    output [63:0] rd_d_0_0;
    output [63:0] rd_d_0_1;
    output [63:0] rd_d_0_2;
    output [63:0] rd_d_0_3;
    output [63:0] rd_d_0_4;
    output [63:0] rd_d_0_5;
    output [63:0] rd_d_0_6;
    output [63:0] rd_d_0_7;
    output [63:0] rd_d_1_0;
    output [63:0] rd_d_1_1;
    output [63:0] rd_d_1_2;
    output [63:0] rd_d_1_3;
    output [63:0] rd_d_1_4;
    output [63:0] rd_d_1_5;
    output [63:0] rd_d_1_6;
    output [63:0] rd_d_1_7;
    output [63:0] rd_d_2_0;
    output [63:0] rd_d_2_1;
    output [63:0] rd_d_2_2;
    output [63:0] rd_d_2_3;
    output [63:0] rd_d_2_4;
    output [63:0] rd_d_2_5;
    output [63:0] rd_d_2_6;
    output [63:0] rd_d_2_7;
    output [63:0] rd_d_3_0;
    output [63:0] rd_d_3_1;
    output [63:0] rd_d_3_2;
    output [63:0] rd_d_3_3;
    output [63:0] rd_d_3_4;
    output [63:0] rd_d_3_5;
    output [63:0] rd_d_3_6;
    output [63:0] rd_d_3_7;

    /* signal declarations */
    wire [63:0] _140;
    wire [63:0] _141;
    wire [63:0] _142;
    wire [63:0] _143;
    wire [63:0] _144;
    wire [63:0] _145;
    wire [63:0] _146;
    wire [5:0] _9;
    wire _134;
    wire [1:0] _135;
    wire [3:0] _136;
    wire [7:0] _137;
    wire [5:0] _11;
    wire _130;
    wire [1:0] _131;
    wire [3:0] _132;
    wire [7:0] _133;
    wire [63:0] _13;
    wire [63:0] _15;
    wire [63:0] _17;
    wire [63:0] _19;
    wire [63:0] _21;
    wire [63:0] _23;
    wire [63:0] _25;
    wire [63:0] _27;
    wire [512:0] _139;
    wire [63:0] _147;
    wire [63:0] _158;
    wire [63:0] _159;
    wire [63:0] _160;
    wire [63:0] _161;
    wire [63:0] _162;
    wire [63:0] _163;
    wire [63:0] _164;
    wire [5:0] _37;
    wire _152;
    wire [1:0] _153;
    wire [3:0] _154;
    wire [7:0] _155;
    wire [5:0] _39;
    wire _148;
    wire [1:0] _149;
    wire [3:0] _150;
    wire [7:0] _151;
    wire [63:0] _41;
    wire [63:0] _43;
    wire [63:0] _45;
    wire [63:0] _47;
    wire [63:0] _49;
    wire [63:0] _51;
    wire [63:0] _53;
    wire [63:0] _55;
    wire [512:0] _157;
    wire [63:0] _165;
    wire [63:0] _176;
    wire [63:0] _177;
    wire [63:0] _178;
    wire [63:0] _179;
    wire [63:0] _180;
    wire [63:0] _181;
    wire [63:0] _182;
    wire [5:0] _65;
    wire _170;
    wire [1:0] _171;
    wire [3:0] _172;
    wire [7:0] _173;
    wire [5:0] _67;
    wire _166;
    wire [1:0] _167;
    wire [3:0] _168;
    wire [7:0] _169;
    wire [63:0] _69;
    wire [63:0] _71;
    wire [63:0] _73;
    wire [63:0] _75;
    wire [63:0] _77;
    wire [63:0] _79;
    wire [63:0] _81;
    wire [63:0] _83;
    wire [512:0] _175;
    wire [63:0] _183;
    wire [63:0] _194;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _197;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _200;
    wire [63:0] _201;
    wire [5:0] _94;
    wire [3:0] _96;
    wire _188;
    wire [1:0] _189;
    wire [3:0] _190;
    wire [7:0] _191;
    wire [5:0] _98;
    wire [3:0] _100;
    wire _184;
    wire [1:0] _185;
    wire [3:0] _186;
    wire [7:0] _187;
    wire [63:0] _102;
    wire [63:0] _104;
    wire [63:0] _106;
    wire [63:0] _108;
    wire [63:0] _110;
    wire [63:0] _112;
    wire [63:0] _114;
    wire [63:0] _116;
    wire _118;
    wire _120;
    wire _122;
    wire _124;
    wire _126;
    wire _128;
    wire [512:0] _193;
    wire _202;

    /* logic */
    assign _140 = _139[512:449];
    assign _141 = _139[448:385];
    assign _142 = _139[384:321];
    assign _143 = _139[320:257];
    assign _144 = _139[256:193];
    assign _145 = _139[192:129];
    assign _146 = _139[128:65];
    assign _9 = rd_addr3;
    assign _134 = _96[3:3];
    assign _135 = { _134, _134 };
    assign _136 = { _135, _135 };
    assign _137 = { _136, _136 };
    assign _11 = wr_addr3;
    assign _130 = _100[3:3];
    assign _131 = { _130, _130 };
    assign _132 = { _131, _131 };
    assign _133 = { _132, _132 };
    assign _13 = wr_d_3_7;
    assign _15 = wr_d_3_6;
    assign _17 = wr_d_3_5;
    assign _19 = wr_d_3_4;
    assign _21 = wr_d_3_3;
    assign _23 = wr_d_3_2;
    assign _25 = wr_d_3_1;
    assign _27 = wr_d_3_0;
    parallel_cores_2
        parallel_cores_2
        ( .clock(_128), .clear(_126), .start(_124), .first_4step_pass(_122), .first_iter(_120), .flip(_118), .wr_d0(_27), .wr_d1(_25), .wr_d2(_23), .wr_d3(_21), .wr_d4(_19), .wr_d5(_17), .wr_d6(_15), .wr_d7(_13), .wr_en(_133), .wr_addr(_11), .rd_en(_137), .rd_addr(_9), .rd_q7(_139[512:449]), .rd_q6(_139[448:385]), .rd_q5(_139[384:321]), .rd_q4(_139[320:257]), .rd_q3(_139[256:193]), .rd_q2(_139[192:129]), .rd_q1(_139[128:65]), .rd_q0(_139[64:1]), .done_(_139[0:0]) );
    assign _147 = _139[64:1];
    assign _158 = _157[512:449];
    assign _159 = _157[448:385];
    assign _160 = _157[384:321];
    assign _161 = _157[320:257];
    assign _162 = _157[256:193];
    assign _163 = _157[192:129];
    assign _164 = _157[128:65];
    assign _37 = rd_addr2;
    assign _152 = _96[2:2];
    assign _153 = { _152, _152 };
    assign _154 = { _153, _153 };
    assign _155 = { _154, _154 };
    assign _39 = wr_addr2;
    assign _148 = _100[2:2];
    assign _149 = { _148, _148 };
    assign _150 = { _149, _149 };
    assign _151 = { _150, _150 };
    assign _41 = wr_d_2_7;
    assign _43 = wr_d_2_6;
    assign _45 = wr_d_2_5;
    assign _47 = wr_d_2_4;
    assign _49 = wr_d_2_3;
    assign _51 = wr_d_2_2;
    assign _53 = wr_d_2_1;
    assign _55 = wr_d_2_0;
    parallel_cores_1
        parallel_cores_1
        ( .clock(_128), .clear(_126), .start(_124), .first_4step_pass(_122), .first_iter(_120), .flip(_118), .wr_d0(_55), .wr_d1(_53), .wr_d2(_51), .wr_d3(_49), .wr_d4(_47), .wr_d5(_45), .wr_d6(_43), .wr_d7(_41), .wr_en(_151), .wr_addr(_39), .rd_en(_155), .rd_addr(_37), .rd_q7(_157[512:449]), .rd_q6(_157[448:385]), .rd_q5(_157[384:321]), .rd_q4(_157[320:257]), .rd_q3(_157[256:193]), .rd_q2(_157[192:129]), .rd_q1(_157[128:65]), .rd_q0(_157[64:1]), .done_(_157[0:0]) );
    assign _165 = _157[64:1];
    assign _176 = _175[512:449];
    assign _177 = _175[448:385];
    assign _178 = _175[384:321];
    assign _179 = _175[320:257];
    assign _180 = _175[256:193];
    assign _181 = _175[192:129];
    assign _182 = _175[128:65];
    assign _65 = rd_addr1;
    assign _170 = _96[1:1];
    assign _171 = { _170, _170 };
    assign _172 = { _171, _171 };
    assign _173 = { _172, _172 };
    assign _67 = wr_addr1;
    assign _166 = _100[1:1];
    assign _167 = { _166, _166 };
    assign _168 = { _167, _167 };
    assign _169 = { _168, _168 };
    assign _69 = wr_d_1_7;
    assign _71 = wr_d_1_6;
    assign _73 = wr_d_1_5;
    assign _75 = wr_d_1_4;
    assign _77 = wr_d_1_3;
    assign _79 = wr_d_1_2;
    assign _81 = wr_d_1_1;
    assign _83 = wr_d_1_0;
    parallel_cores_0
        parallel_cores_0
        ( .clock(_128), .clear(_126), .start(_124), .first_4step_pass(_122), .first_iter(_120), .flip(_118), .wr_d0(_83), .wr_d1(_81), .wr_d2(_79), .wr_d3(_77), .wr_d4(_75), .wr_d5(_73), .wr_d6(_71), .wr_d7(_69), .wr_en(_169), .wr_addr(_67), .rd_en(_173), .rd_addr(_65), .rd_q7(_175[512:449]), .rd_q6(_175[448:385]), .rd_q5(_175[384:321]), .rd_q4(_175[320:257]), .rd_q3(_175[256:193]), .rd_q2(_175[192:129]), .rd_q1(_175[128:65]), .rd_q0(_175[64:1]), .done_(_175[0:0]) );
    assign _183 = _175[64:1];
    assign _194 = _193[512:449];
    assign _195 = _193[448:385];
    assign _196 = _193[384:321];
    assign _197 = _193[320:257];
    assign _198 = _193[256:193];
    assign _199 = _193[192:129];
    assign _200 = _193[128:65];
    assign _201 = _193[64:1];
    assign _94 = rd_addr0;
    assign _96 = rd_en;
    assign _188 = _96[0:0];
    assign _189 = { _188, _188 };
    assign _190 = { _189, _189 };
    assign _191 = { _190, _190 };
    assign _98 = wr_addr0;
    assign _100 = wr_en;
    assign _184 = _100[0:0];
    assign _185 = { _184, _184 };
    assign _186 = { _185, _185 };
    assign _187 = { _186, _186 };
    assign _102 = wr_d_0_7;
    assign _104 = wr_d_0_6;
    assign _106 = wr_d_0_5;
    assign _108 = wr_d_0_4;
    assign _110 = wr_d_0_3;
    assign _112 = wr_d_0_2;
    assign _114 = wr_d_0_1;
    assign _116 = wr_d_0_0;
    assign _118 = flip;
    assign _120 = first_iter;
    assign _122 = first_4step_pass;
    assign _124 = start;
    assign _126 = clear;
    assign _128 = clock;
    parallel_cores
        parallel_cores
        ( .clock(_128), .clear(_126), .start(_124), .first_4step_pass(_122), .first_iter(_120), .flip(_118), .wr_d0(_116), .wr_d1(_114), .wr_d2(_112), .wr_d3(_110), .wr_d4(_108), .wr_d5(_106), .wr_d6(_104), .wr_d7(_102), .wr_en(_187), .wr_addr(_98), .rd_en(_191), .rd_addr(_94), .rd_q7(_193[512:449]), .rd_q6(_193[448:385]), .rd_q5(_193[384:321]), .rd_q4(_193[320:257]), .rd_q3(_193[256:193]), .rd_q2(_193[192:129]), .rd_q1(_193[128:65]), .rd_q0(_193[64:1]), .done_(_193[0:0]) );
    assign _202 = _193[0:0];

    /* aliases */

    /* output assignments */
    assign done_ = _202;
    assign rd_d_0_0 = _201;
    assign rd_d_0_1 = _200;
    assign rd_d_0_2 = _199;
    assign rd_d_0_3 = _198;
    assign rd_d_0_4 = _197;
    assign rd_d_0_5 = _196;
    assign rd_d_0_6 = _195;
    assign rd_d_0_7 = _194;
    assign rd_d_1_0 = _183;
    assign rd_d_1_1 = _182;
    assign rd_d_1_2 = _181;
    assign rd_d_1_3 = _180;
    assign rd_d_1_4 = _179;
    assign rd_d_1_5 = _178;
    assign rd_d_1_6 = _177;
    assign rd_d_1_7 = _176;
    assign rd_d_2_0 = _165;
    assign rd_d_2_1 = _164;
    assign rd_d_2_2 = _163;
    assign rd_d_2_3 = _162;
    assign rd_d_2_4 = _161;
    assign rd_d_2_5 = _160;
    assign rd_d_2_6 = _159;
    assign rd_d_2_7 = _158;
    assign rd_d_3_0 = _147;
    assign rd_d_3_1 = _146;
    assign rd_d_3_2 = _145;
    assign rd_d_3_3 = _144;
    assign rd_d_3_4 = _143;
    assign rd_d_3_5 = _142;
    assign rd_d_3_6 = _141;
    assign rd_d_3_7 = _140;

endmodule
module kernel (
    data_in_tdata,
    data_in_tvalid,
    first_4step_pass,
    start,
    data_out_dest_tready,
    clear,
    clock,
    data_in_tkeep,
    data_in_tlast,
    data_in_tstrb,
    data_out_tvalid,
    data_out_tdata,
    data_out_tkeep,
    data_out_tstrb,
    data_out_tlast,
    data_in_dest_tready,
    done_
);

    input [511:0] data_in_tdata;
    input data_in_tvalid;
    input first_4step_pass;
    input start;
    input data_out_dest_tready;
    input clear;
    input clock;
    input [63:0] data_in_tkeep;
    input data_in_tlast;
    input [63:0] data_in_tstrb;
    output data_out_tvalid;
    output [511:0] data_out_tdata;
    output [63:0] data_out_tkeep;
    output [63:0] data_out_tstrb;
    output data_out_tlast;
    output data_in_dest_tready;
    output done_;

    /* signal declarations */
    wire _33;
    wire _34;
    wire gnd = 1'b0;
    wire [63:0] _36 = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    wire [63:0] _37 = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    wire [511:0] _245 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _244 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _242 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _241 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _238 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _237 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _235 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _234 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _232 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _231 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _229;
    wire [63:0] _228;
    wire [63:0] _227;
    wire [63:0] _226;
    wire [63:0] _225;
    wire [63:0] _224;
    wire [63:0] _223;
    wire [63:0] _222;
    wire [511:0] _230;
    (* keep="TRUE" *)
    reg [511:0] _233;
    (* keep="TRUE" *)
    reg [511:0] _236;
    (* keep="TRUE" *)
    reg [511:0] _239;
    wire [511:0] _220 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _219 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _217 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _216 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _214 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _213 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _211;
    wire [63:0] _210;
    wire [63:0] _209;
    wire [63:0] _208;
    wire [63:0] _207;
    wire [63:0] _206;
    wire [63:0] _205;
    wire [63:0] _204;
    wire [511:0] _212;
    (* keep="TRUE" *)
    reg [511:0] _215;
    (* keep="TRUE" *)
    reg [511:0] _218;
    (* keep="TRUE" *)
    reg [511:0] _221;
    wire [511:0] _202 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _201 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _199 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _198 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _196 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _195 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _193;
    wire [63:0] _192;
    wire [63:0] _191;
    wire [63:0] _190;
    wire [63:0] _189;
    wire [63:0] _188;
    wire [63:0] _187;
    wire [63:0] _186;
    wire [511:0] _194;
    (* keep="TRUE" *)
    reg [511:0] _197;
    (* keep="TRUE" *)
    reg [511:0] _200;
    (* keep="TRUE" *)
    reg [511:0] _203;
    wire [511:0] _184 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _183 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _181 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _180 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _178 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _177 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _175;
    wire [63:0] _174;
    wire [63:0] _173;
    wire [63:0] _172;
    wire [63:0] _171;
    wire [63:0] _170;
    wire [63:0] _169;
    wire [63:0] _168;
    wire [511:0] _176;
    (* keep="TRUE" *)
    reg [511:0] _179;
    (* keep="TRUE" *)
    reg [511:0] _182;
    (* keep="TRUE" *)
    reg [511:0] _185;
    wire [1:0] _62 = 2'b00;
    wire [1:0] _61 = 2'b00;
    wire [1:0] _59 = 2'b00;
    wire [1:0] _58 = 2'b00;
    wire [1:0] _56 = 2'b00;
    wire [1:0] _55 = 2'b00;
    wire [1:0] _53 = 2'b00;
    wire [1:0] _52 = 2'b00;
    wire [1:0] _50 = 2'b00;
    wire [1:0] _49 = 2'b00;
    wire [1:0] _47 = 2'b00;
    wire [1:0] _46 = 2'b00;
    wire [3:0] _42 = 4'b0000;
    wire _43;
    wire _44;
    wire [1:0] _40 = 2'b00;
    wire [1:0] _39 = 2'b00;
    wire [1:0] _38;
    reg [1:0] _45;
    reg [1:0] _48;
    reg [1:0] _51;
    reg [1:0] _54;
    reg [1:0] _57;
    reg [1:0] _60;
    reg [1:0] _63;
    reg [511:0] _240;
    reg [511:0] _243;
    reg [511:0] _246;
    wire [5:0] _164 = 6'b000000;
    wire [5:0] _163 = 6'b000000;
    wire [5:0] _161 = 6'b000000;
    wire [5:0] _160 = 6'b000000;
    wire [5:0] _158 = 6'b000000;
    wire [5:0] _157 = 6'b000000;
    (* keep="TRUE" *)
    reg [5:0] _159;
    (* keep="TRUE" *)
    reg [5:0] _162;
    (* keep="TRUE" *)
    reg [5:0] _165;
    wire [5:0] _155 = 6'b000000;
    wire [5:0] _154 = 6'b000000;
    wire [5:0] _152 = 6'b000000;
    wire [5:0] _151 = 6'b000000;
    wire [5:0] _149 = 6'b000000;
    wire [5:0] _148 = 6'b000000;
    (* keep="TRUE" *)
    reg [5:0] _150;
    (* keep="TRUE" *)
    reg [5:0] _153;
    (* keep="TRUE" *)
    reg [5:0] _156;
    wire [5:0] _146 = 6'b000000;
    wire [5:0] _145 = 6'b000000;
    wire [5:0] _143 = 6'b000000;
    wire [5:0] _142 = 6'b000000;
    wire [5:0] _140 = 6'b000000;
    wire [5:0] _139 = 6'b000000;
    (* keep="TRUE" *)
    reg [5:0] _141;
    (* keep="TRUE" *)
    reg [5:0] _144;
    (* keep="TRUE" *)
    reg [5:0] _147;
    wire [5:0] _137 = 6'b000000;
    wire [5:0] _136 = 6'b000000;
    wire [5:0] _134 = 6'b000000;
    wire [5:0] _133 = 6'b000000;
    wire [5:0] _131 = 6'b000000;
    wire [5:0] _130 = 6'b000000;
    wire [5:0] _129;
    (* keep="TRUE" *)
    reg [5:0] _132;
    (* keep="TRUE" *)
    reg [5:0] _135;
    (* keep="TRUE" *)
    reg [5:0] _138;
    wire [3:0] _127 = 4'b0000;
    wire [3:0] _126 = 4'b0000;
    wire [3:0] _124 = 4'b0000;
    wire [3:0] _123 = 4'b0000;
    wire [3:0] _121 = 4'b0000;
    wire [3:0] _120 = 4'b0000;
    wire [3:0] _41;
    (* keep="TRUE" *)
    reg [3:0] _122;
    (* keep="TRUE" *)
    reg [3:0] _125;
    (* keep="TRUE" *)
    reg [3:0] _128;
    wire [5:0] _118 = 6'b000000;
    wire [5:0] _117 = 6'b000000;
    wire [5:0] _115 = 6'b000000;
    wire [5:0] _114 = 6'b000000;
    (* keep="TRUE" *)
    reg [5:0] _116;
    (* keep="TRUE" *)
    reg [5:0] _119;
    wire [5:0] _112 = 6'b000000;
    wire [5:0] _111 = 6'b000000;
    wire [5:0] _109 = 6'b000000;
    wire [5:0] _108 = 6'b000000;
    (* keep="TRUE" *)
    reg [5:0] _110;
    (* keep="TRUE" *)
    reg [5:0] _113;
    wire [5:0] _106 = 6'b000000;
    wire [5:0] _105 = 6'b000000;
    wire [5:0] _103 = 6'b000000;
    wire [5:0] _102 = 6'b000000;
    (* keep="TRUE" *)
    reg [5:0] _104;
    (* keep="TRUE" *)
    reg [5:0] _107;
    wire [5:0] _100 = 6'b000000;
    wire [5:0] _99 = 6'b000000;
    wire [5:0] _97 = 6'b000000;
    wire [5:0] _96 = 6'b000000;
    wire [5:0] _95;
    (* keep="TRUE" *)
    reg [5:0] _98;
    (* keep="TRUE" *)
    reg [5:0] _101;
    wire [3:0] _93 = 4'b0000;
    wire [3:0] _92 = 4'b0000;
    wire [3:0] _90 = 4'b0000;
    wire [3:0] _89 = 4'b0000;
    wire [3:0] _88;
    (* keep="TRUE" *)
    reg [3:0] _91;
    (* keep="TRUE" *)
    reg [3:0] _94;
    wire [63:0] _87;
    wire [127:0] _85;
    wire [63:0] _86;
    wire [191:0] _83;
    wire [63:0] _84;
    wire [255:0] _81;
    wire [63:0] _82;
    wire [319:0] _79;
    wire [63:0] _80;
    wire [383:0] _77;
    wire [63:0] _78;
    wire [447:0] _75;
    wire [63:0] _76;
    wire [511:0] _72 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _71 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [511:0] _68 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _67 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _8;
    reg [511:0] _70;
    reg [511:0] _73;
    wire [63:0] _74;
    wire _66;
    wire _65;
    wire _64;
    wire [2048:0] _167;
    wire _247;
    wire _9;
    wire _30;
    wire _248;
    wire _10;
    wire _12;
    wire _14;
    wire [11:0] _26;
    wire _27;
    wire _16;
    wire [5:0] _32;
    wire _249;
    wire _17;
    wire _19;
    wire _21;
    wire _23;
    wire [13:0] _29;
    wire _250;

    /* logic */
    assign _33 = _32[0:0];
    assign _34 = _26[1:1];
    assign _229 = _167[1600:1537];
    assign _228 = _167[1664:1601];
    assign _227 = _167[1728:1665];
    assign _226 = _167[1792:1729];
    assign _225 = _167[1856:1793];
    assign _224 = _167[1920:1857];
    assign _223 = _167[1984:1921];
    assign _222 = _167[2048:1985];
    assign _230 = { _222, _223, _224, _225, _226, _227, _228, _229 };
    always @(posedge _23) begin
        if (_44)
            _233 <= _230;
    end
    always @(posedge _23) begin
        if (_44)
            _236 <= _233;
    end
    always @(posedge _23) begin
        if (_44)
            _239 <= _236;
    end
    assign _211 = _167[1088:1025];
    assign _210 = _167[1152:1089];
    assign _209 = _167[1216:1153];
    assign _208 = _167[1280:1217];
    assign _207 = _167[1344:1281];
    assign _206 = _167[1408:1345];
    assign _205 = _167[1472:1409];
    assign _204 = _167[1536:1473];
    assign _212 = { _204, _205, _206, _207, _208, _209, _210, _211 };
    always @(posedge _23) begin
        if (_44)
            _215 <= _212;
    end
    always @(posedge _23) begin
        if (_44)
            _218 <= _215;
    end
    always @(posedge _23) begin
        if (_44)
            _221 <= _218;
    end
    assign _193 = _167[576:513];
    assign _192 = _167[640:577];
    assign _191 = _167[704:641];
    assign _190 = _167[768:705];
    assign _189 = _167[832:769];
    assign _188 = _167[896:833];
    assign _187 = _167[960:897];
    assign _186 = _167[1024:961];
    assign _194 = { _186, _187, _188, _189, _190, _191, _192, _193 };
    always @(posedge _23) begin
        if (_44)
            _197 <= _194;
    end
    always @(posedge _23) begin
        if (_44)
            _200 <= _197;
    end
    always @(posedge _23) begin
        if (_44)
            _203 <= _200;
    end
    assign _175 = _167[64:1];
    assign _174 = _167[128:65];
    assign _173 = _167[192:129];
    assign _172 = _167[256:193];
    assign _171 = _167[320:257];
    assign _170 = _167[384:321];
    assign _169 = _167[448:385];
    assign _168 = _167[512:449];
    assign _176 = { _168, _169, _170, _171, _172, _173, _174, _175 };
    always @(posedge _23) begin
        if (_44)
            _179 <= _176;
    end
    always @(posedge _23) begin
        if (_44)
            _182 <= _179;
    end
    always @(posedge _23) begin
        if (_44)
            _185 <= _182;
    end
    assign _43 = _41 == _42;
    assign _44 = ~ _43;
    assign _38 = _29[13:12];
    always @(posedge _23) begin
        if (_44)
            _45 <= _38;
    end
    always @(posedge _23) begin
        if (_44)
            _48 <= _45;
    end
    always @(posedge _23) begin
        if (_44)
            _51 <= _48;
    end
    always @(posedge _23) begin
        if (_44)
            _54 <= _51;
    end
    always @(posedge _23) begin
        if (_44)
            _57 <= _54;
    end
    always @(posedge _23) begin
        if (_44)
            _60 <= _57;
    end
    always @(posedge _23) begin
        if (_44)
            _63 <= _60;
    end
    always @* begin
        case (_63)
        0: _240 <= _185;
        1: _240 <= _203;
        2: _240 <= _221;
        default: _240 <= _239;
        endcase
    end
    always @(posedge _23) begin
        if (_44)
            _243 <= _240;
    end
    always @(posedge _23) begin
        if (_44)
            _246 <= _243;
    end
    always @(posedge _23) begin
        _159 <= _129;
    end
    always @(posedge _23) begin
        _162 <= _159;
    end
    always @(posedge _23) begin
        _165 <= _162;
    end
    always @(posedge _23) begin
        _150 <= _129;
    end
    always @(posedge _23) begin
        _153 <= _150;
    end
    always @(posedge _23) begin
        _156 <= _153;
    end
    always @(posedge _23) begin
        _141 <= _129;
    end
    always @(posedge _23) begin
        _144 <= _141;
    end
    always @(posedge _23) begin
        _147 <= _144;
    end
    assign _129 = _29[7:2];
    always @(posedge _23) begin
        _132 <= _129;
    end
    always @(posedge _23) begin
        _135 <= _132;
    end
    always @(posedge _23) begin
        _138 <= _135;
    end
    assign _41 = _29[11:8];
    always @(posedge _23) begin
        _122 <= _41;
    end
    always @(posedge _23) begin
        _125 <= _122;
    end
    always @(posedge _23) begin
        _128 <= _125;
    end
    always @(posedge _23) begin
        _116 <= _95;
    end
    always @(posedge _23) begin
        _119 <= _116;
    end
    always @(posedge _23) begin
        _110 <= _95;
    end
    always @(posedge _23) begin
        _113 <= _110;
    end
    always @(posedge _23) begin
        _104 <= _95;
    end
    always @(posedge _23) begin
        _107 <= _104;
    end
    assign _95 = _26[7:2];
    always @(posedge _23) begin
        _98 <= _95;
    end
    always @(posedge _23) begin
        _101 <= _98;
    end
    assign _88 = _26[11:8];
    always @(posedge _23) begin
        _91 <= _88;
    end
    always @(posedge _23) begin
        _94 <= _91;
    end
    assign _87 = _85[127:64];
    assign _85 = _83[191:64];
    assign _86 = _85[63:0];
    assign _83 = _81[255:64];
    assign _84 = _83[63:0];
    assign _81 = _79[319:64];
    assign _82 = _81[63:0];
    assign _79 = _77[383:64];
    assign _80 = _79[63:0];
    assign _77 = _75[447:64];
    assign _78 = _77[63:0];
    assign _75 = _73[511:64];
    assign _76 = _75[63:0];
    assign _8 = data_in_tdata;
    always @(posedge _23) begin
        _70 <= _8;
    end
    always @(posedge _23) begin
        _73 <= _70;
    end
    assign _74 = _73[63:0];
    assign _66 = _32[5:5];
    assign _65 = _32[4:4];
    assign _64 = _32[3:3];
    multi_parallel_cores
        multi_parallel_cores
        ( .clock(_23), .clear(_21), .start(_64), .first_4step_pass(_14), .first_iter(_65), .flip(_66), .wr_d_0_0(_74), .wr_d_0_1(_76), .wr_d_0_2(_78), .wr_d_0_3(_80), .wr_d_0_4(_82), .wr_d_0_5(_84), .wr_d_0_6(_86), .wr_d_0_7(_87), .wr_d_1_0(_74), .wr_d_1_1(_76), .wr_d_1_2(_78), .wr_d_1_3(_80), .wr_d_1_4(_82), .wr_d_1_5(_84), .wr_d_1_6(_86), .wr_d_1_7(_87), .wr_d_2_0(_74), .wr_d_2_1(_76), .wr_d_2_2(_78), .wr_d_2_3(_80), .wr_d_2_4(_82), .wr_d_2_5(_84), .wr_d_2_6(_86), .wr_d_2_7(_87), .wr_d_3_0(_74), .wr_d_3_1(_76), .wr_d_3_2(_78), .wr_d_3_3(_80), .wr_d_3_4(_82), .wr_d_3_5(_84), .wr_d_3_6(_86), .wr_d_3_7(_87), .wr_en(_94), .wr_addr0(_101), .wr_addr1(_107), .wr_addr2(_113), .wr_addr3(_119), .rd_en(_128), .rd_addr0(_138), .rd_addr1(_147), .rd_addr2(_156), .rd_addr3(_165), .rd_d_3_7(_167[2048:1985]), .rd_d_3_6(_167[1984:1921]), .rd_d_3_5(_167[1920:1857]), .rd_d_3_4(_167[1856:1793]), .rd_d_3_3(_167[1792:1729]), .rd_d_3_2(_167[1728:1665]), .rd_d_3_1(_167[1664:1601]), .rd_d_3_0(_167[1600:1537]), .rd_d_2_7(_167[1536:1473]), .rd_d_2_6(_167[1472:1409]), .rd_d_2_5(_167[1408:1345]), .rd_d_2_4(_167[1344:1281]), .rd_d_2_3(_167[1280:1217]), .rd_d_2_2(_167[1216:1153]), .rd_d_2_1(_167[1152:1089]), .rd_d_2_0(_167[1088:1025]), .rd_d_1_7(_167[1024:961]), .rd_d_1_6(_167[960:897]), .rd_d_1_5(_167[896:833]), .rd_d_1_4(_167[832:769]), .rd_d_1_3(_167[768:705]), .rd_d_1_2(_167[704:641]), .rd_d_1_1(_167[640:577]), .rd_d_1_0(_167[576:513]), .rd_d_0_7(_167[512:449]), .rd_d_0_6(_167[448:385]), .rd_d_0_5(_167[384:321]), .rd_d_0_4(_167[320:257]), .rd_d_0_3(_167[256:193]), .rd_d_0_2(_167[192:129]), .rd_d_0_1(_167[128:65]), .rd_d_0_0(_167[64:1]), .done_(_167[0:0]) );
    assign _247 = _167[0:0];
    assign _9 = _247;
    assign _30 = _29[0:0];
    assign _248 = _32[1:1];
    assign _10 = _248;
    assign _12 = data_in_tvalid;
    assign _14 = first_4step_pass;
    load_sm
        load_sm
        ( .clock(_23), .clear(_21), .first_4step_pass(_14), .tvalid(_12), .start(_10), .wr_en(_26[11:8]), .wr_addr(_26[7:2]), .tready(_26[1:1]), .done_(_26[0:0]) );
    assign _27 = _26[0:0];
    assign _16 = start;
    controller
        controller
        ( .clock(_23), .clear(_21), .start(_16), .input_done(_27), .output_done(_30), .cores_done(_9), .flip(_32[5:5]), .first_iter(_32[4:4]), .start_cores(_32[3:3]), .start_output(_32[2:2]), .start_input(_32[1:1]), .done_(_32[0:0]) );
    assign _249 = _32[2:2];
    assign _17 = _249;
    assign _19 = data_out_dest_tready;
    assign _21 = clear;
    assign _23 = clock;
    store_sm
        store_sm
        ( .clock(_23), .clear(_21), .tready(_19), .start(_17), .block(_29[13:12]), .rd_en(_29[11:8]), .rd_addr(_29[7:2]), .tvalid(_29[1:1]), .done_(_29[0:0]) );
    assign _250 = _29[1:1];

    /* aliases */

    /* output assignments */
    assign data_out_tvalid = _250;
    assign data_out_tdata = _246;
    assign data_out_tkeep = _37;
    assign data_out_tstrb = _36;
    assign data_out_tlast = gnd;
    assign data_in_dest_tready = _34;
    assign done_ = _33;

endmodule
module transposer_memories (
    write_enable,
    write_data,
    write_address,
    clock,
    read_address,
    read_data0,
    read_data1,
    read_data2,
    read_data3,
    read_data4,
    read_data5,
    read_data6,
    read_data7
);

    input [7:0] write_enable;
    input [511:0] write_data;
    input [2:0] write_address;
    input clock;
    input [2:0] read_address;
    (* RAM_STYLE="distributed" *)
    output [511:0] read_data0;
    (* RAM_STYLE="distributed" *)
    output [511:0] read_data1;
    (* RAM_STYLE="distributed" *)
    output [511:0] read_data2;
    (* RAM_STYLE="distributed" *)
    output [511:0] read_data3;
    (* RAM_STYLE="distributed" *)
    output [511:0] read_data4;
    (* RAM_STYLE="distributed" *)
    output [511:0] read_data5;
    (* RAM_STYLE="distributed" *)
    output [511:0] read_data6;
    (* RAM_STYLE="distributed" *)
    output [511:0] read_data7;

    /* signal declarations */
    wire _19;
    reg [511:0] _20[0:7];
    wire [511:0] _21;
    wire _22;
    reg [511:0] _23[0:7];
    wire [511:0] _24;
    wire _25;
    reg [511:0] _26[0:7];
    wire [511:0] _27;
    wire _28;
    reg [511:0] _29[0:7];
    wire [511:0] _30;
    wire _31;
    reg [511:0] _32[0:7];
    wire [511:0] _33;
    wire _34;
    reg [511:0] _35[0:7];
    wire [511:0] _36;
    wire _37;
    reg [511:0] _38[0:7];
    wire [511:0] _39;
    wire [7:0] _9;
    wire _40;
    wire [511:0] _11;
    wire [2:0] _13;
    wire _15;
    reg [511:0] _41[0:7];
    wire [2:0] _17;
    wire [511:0] _42;

    /* logic */
    assign _19 = _9[7:7];
    always @(posedge _15) begin
        if (_19)
            _20[_13] <= _11;
    end
    assign _21 = _20[_17];
    assign _22 = _9[6:6];
    always @(posedge _15) begin
        if (_22)
            _23[_13] <= _11;
    end
    assign _24 = _23[_17];
    assign _25 = _9[5:5];
    always @(posedge _15) begin
        if (_25)
            _26[_13] <= _11;
    end
    assign _27 = _26[_17];
    assign _28 = _9[4:4];
    always @(posedge _15) begin
        if (_28)
            _29[_13] <= _11;
    end
    assign _30 = _29[_17];
    assign _31 = _9[3:3];
    always @(posedge _15) begin
        if (_31)
            _32[_13] <= _11;
    end
    assign _33 = _32[_17];
    assign _34 = _9[2:2];
    always @(posedge _15) begin
        if (_34)
            _35[_13] <= _11;
    end
    assign _36 = _35[_17];
    assign _37 = _9[1:1];
    always @(posedge _15) begin
        if (_37)
            _38[_13] <= _11;
    end
    assign _39 = _38[_17];
    assign _9 = write_enable;
    assign _40 = _9[0:0];
    assign _11 = write_data;
    assign _13 = write_address;
    assign _15 = clock;
    always @(posedge _15) begin
        if (_40)
            _41[_13] <= _11;
    end
    assign _17 = read_address;
    assign _42 = _41[_17];

    /* aliases */

    /* output assignments */
    assign read_data0 = _42;
    assign read_data1 = _39;
    assign read_data2 = _36;
    assign read_data3 = _33;
    assign read_data4 = _30;
    assign read_data5 = _27;
    assign read_data6 = _24;
    assign read_data7 = _21;

endmodule
module transposer (
    in_tdata,
    in_tvalid,
    clear,
    clock,
    out_tready,
    in_tkeep,
    in_tlast,
    in_tstrb,
    out_tvalid,
    out_tdata,
    out_tkeep,
    out_tstrb,
    out_tlast,
    in_tready
);

    input [511:0] in_tdata;
    input in_tvalid;
    input clear;
    input clock;
    input out_tready;
    input [63:0] in_tkeep;
    input in_tlast;
    input [63:0] in_tstrb;
    output out_tvalid;
    output [511:0] out_tdata;
    output [63:0] out_tkeep;
    output [63:0] out_tstrb;
    output out_tlast;
    output in_tready;

    /* signal declarations */
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    wire _72 = 1'b1;
    wire _73;
    wire _59 = 1'b0;
    wire _60;
    wire _61;
    wire _62;
    wire _46;
    wire _63;
    wire _44;
    wire _74;
    wire _1;
    reg _49;
    wire _2;
    wire gnd = 1'b0;
    wire _4;
    wire [63:0] _76 = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    wire [63:0] _6;
    wire [63:0] _77 = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    wire [63:0] _8;
    wire [63:0] _225;
    wire [127:0] _223;
    wire [63:0] _224;
    wire [191:0] _221;
    wire [63:0] _222;
    wire [255:0] _219;
    wire [63:0] _220;
    wire [319:0] _217;
    wire [63:0] _218;
    wire [383:0] _215;
    wire [63:0] _216;
    wire [447:0] _213;
    wire [63:0] _214;
    wire [511:0] _211;
    wire [63:0] _212;
    reg [63:0] _226;
    wire [63:0] _209;
    wire [127:0] _207;
    wire [63:0] _208;
    wire [191:0] _205;
    wire [63:0] _206;
    wire [255:0] _203;
    wire [63:0] _204;
    wire [319:0] _201;
    wire [63:0] _202;
    wire [383:0] _199;
    wire [63:0] _200;
    wire [447:0] _197;
    wire [63:0] _198;
    wire [511:0] _195;
    wire [63:0] _196;
    reg [63:0] _210;
    wire [63:0] _193;
    wire [127:0] _191;
    wire [63:0] _192;
    wire [191:0] _189;
    wire [63:0] _190;
    wire [255:0] _187;
    wire [63:0] _188;
    wire [319:0] _185;
    wire [63:0] _186;
    wire [383:0] _183;
    wire [63:0] _184;
    wire [447:0] _181;
    wire [63:0] _182;
    wire [511:0] _179;
    wire [63:0] _180;
    reg [63:0] _194;
    wire [63:0] _177;
    wire [127:0] _175;
    wire [63:0] _176;
    wire [191:0] _173;
    wire [63:0] _174;
    wire [255:0] _171;
    wire [63:0] _172;
    wire [319:0] _169;
    wire [63:0] _170;
    wire [383:0] _167;
    wire [63:0] _168;
    wire [447:0] _165;
    wire [63:0] _166;
    wire [511:0] _163;
    wire [63:0] _164;
    reg [63:0] _178;
    wire [63:0] _161;
    wire [127:0] _159;
    wire [63:0] _160;
    wire [191:0] _157;
    wire [63:0] _158;
    wire [255:0] _155;
    wire [63:0] _156;
    wire [319:0] _153;
    wire [63:0] _154;
    wire [383:0] _151;
    wire [63:0] _152;
    wire [447:0] _149;
    wire [63:0] _150;
    wire [511:0] _147;
    wire [63:0] _148;
    reg [63:0] _162;
    wire [63:0] _145;
    wire [127:0] _143;
    wire [63:0] _144;
    wire [191:0] _141;
    wire [63:0] _142;
    wire [255:0] _139;
    wire [63:0] _140;
    wire [319:0] _137;
    wire [63:0] _138;
    wire [383:0] _135;
    wire [63:0] _136;
    wire [447:0] _133;
    wire [63:0] _134;
    wire [511:0] _131;
    wire [63:0] _132;
    reg [63:0] _146;
    wire [63:0] _129;
    wire [127:0] _127;
    wire [63:0] _128;
    wire [191:0] _125;
    wire [63:0] _126;
    wire [255:0] _123;
    wire [63:0] _124;
    wire [319:0] _121;
    wire [63:0] _122;
    wire [383:0] _119;
    wire [63:0] _120;
    wire [447:0] _117;
    wire [63:0] _118;
    wire [511:0] _115;
    wire [63:0] _116;
    reg [63:0] _130;
    wire [63:0] _113;
    wire [127:0] _111;
    wire [63:0] _112;
    wire [191:0] _109;
    wire [63:0] _110;
    wire [255:0] _107;
    wire [63:0] _108;
    wire [319:0] _105;
    wire [63:0] _106;
    wire [383:0] _103;
    wire [63:0] _104;
    wire [447:0] _101;
    wire [63:0] _102;
    wire [511:0] _11;
    wire [511:0] _12;
    wire _78;
    wire _79;
    wire [1:0] _80;
    wire [3:0] _81;
    wire [7:0] _82;
    wire [7:0] _83;
    wire [7:0] _13;
    wire _84;
    wire [2:0] _85;
    wire [2:0] _14;
    wire _89;
    wire [2:0] _93;
    wire [2:0] _15;
    wire [4095:0] _98;
    wire [511:0] _99;
    wire [63:0] _100;
    reg [63:0] _114;
    wire [511:0] _227;
    wire [511:0] _16;
    wire _314 = 1'b0;
    wire _313 = 1'b0;
    wire _321 = 1'b1;
    wire _322;
    wire _316 = 1'b0;
    wire _317;
    wire _318;
    wire _319;
    wire _312;
    wire _320;
    wire _265 = 1'b0;
    wire _264 = 1'b0;
    wire [1:0] _305 = 2'b10;
    wire [1:0] _306;
    wire _307;
    wire [1:0] _302 = 2'b01;
    wire [1:0] _65 = 2'b00;
    wire [1:0] _64 = 2'b00;
    wire [1:0] _258 = 2'b01;
    wire [1:0] _259;
    wire [1:0] _260;
    wire [1:0] _261;
    wire [1:0] _262;
    wire _40 = 1'b0;
    wire _39 = 1'b0;
    wire _255;
    wire [7:0] _56 = 8'b00000000;
    wire [7:0] _55 = 8'b00000000;
    wire [7:0] _239 = 8'b00000001;
    wire [7:0] _238 = 8'b00000000;
    wire [1:0] _68 = 2'b01;
    wire [1:0] _69;
    wire _70;
    wire [1:0] rd_pos;
    wire _67;
    wire _71;
    wire [7:0] _240;
    wire [7:0] _233 = 8'b00000000;
    wire _231 = 1'b0;
    wire [6:0] _230;
    wire [7:0] _232;
    wire [7:0] _234;
    wire [7:0] _235;
    wire [7:0] _236;
    wire _229;
    wire [7:0] _237;
    wire _228;
    wire [7:0] _241;
    wire [7:0] _19;
    reg [7:0] _57;
    wire _58;
    wire _251;
    wire [1:0] _53 = 2'b11;
    wire [1:0] _51 = 2'b00;
    wire [1:0] _50 = 2'b00;
    wire [1:0] _245 = 2'b00;
    wire [1:0] _243 = 2'b01;
    wire [1:0] _244;
    wire [1:0] _246;
    wire [1:0] _247;
    wire _242;
    wire [1:0] _248;
    wire [1:0] _20;
    reg [1:0] _52;
    wire _54;
    wire _252;
    wire _22;
    wire _253;
    wire _45 = 1'b1;
    wire _250;
    wire _254;
    wire _43 = 1'b0;
    wire _249;
    wire _256;
    wire _23;
    reg _42;
    wire _257;
    wire [1:0] _263;
    wire [1:0] _24;
    reg [1:0] _66;
    wire [1:0] wr_pos;
    wire [1:0] _303;
    wire [1:0] _87 = 2'b00;
    wire [1:0] _86 = 2'b00;
    wire [1:0] _273 = 2'b01;
    wire [1:0] _274;
    wire [1:0] _275;
    wire [1:0] _276;
    wire [1:0] _277;
    wire _268;
    wire [1:0] _278;
    wire [1:0] _26;
    reg [1:0] _88;
    wire _304;
    wire _308;
    wire _309;
    wire [1:0] _271 = 2'b11;
    wire [1:0] _91 = 2'b00;
    wire [1:0] _90 = 2'b00;
    wire [1:0] _289 = 2'b00;
    wire [1:0] _284 = 2'b00;
    wire [1:0] _282 = 2'b01;
    wire [1:0] _283;
    wire [1:0] _285;
    wire [1:0] _286;
    wire [1:0] _287;
    wire _281;
    wire [1:0] _288;
    wire _280;
    wire [1:0] _290;
    wire [1:0] _27;
    reg [1:0] _92;
    wire _272;
    wire _298;
    wire [2:0] _269 = 3'b111;
    wire vdd = 1'b1;
    wire [2:0] _95 = 3'b000;
    wire _29;
    wire [2:0] _94 = 3'b000;
    wire _31;
    wire [2:0] _292 = 3'b001;
    wire [2:0] _293;
    wire [2:0] _294;
    wire _291;
    wire [2:0] _295;
    wire [2:0] _32;
    reg [2:0] element_offset;
    wire _270;
    wire _299;
    wire _34;
    wire _300;
    wire _267 = 1'b1;
    wire _297;
    wire _301;
    wire _279 = 1'b0;
    wire _296;
    wire _310;
    wire _35;
    reg _266;
    wire _311;
    wire _323;
    wire _36;
    reg _315;
    wire _37;

    /* logic */
    assign _73 = _71 ? _72 : _49;
    assign _60 = _58 ? _59 : _49;
    assign _61 = _54 ? _60 : _49;
    assign _62 = _22 ? _61 : _49;
    assign _46 = _42 == _45;
    assign _63 = _46 ? _62 : _49;
    assign _44 = _42 == _43;
    assign _74 = _44 ? _73 : _63;
    assign _1 = _74;
    always @(posedge _31) begin
        if (_29)
            _49 <= _48;
        else
            _49 <= _1;
    end
    assign _2 = _49;
    assign _4 = gnd;
    assign _6 = _76;
    assign _8 = _77;
    assign _225 = _223[127:64];
    assign _223 = _221[191:64];
    assign _224 = _223[63:0];
    assign _221 = _219[255:64];
    assign _222 = _221[63:0];
    assign _219 = _217[319:64];
    assign _220 = _219[63:0];
    assign _217 = _215[383:64];
    assign _218 = _217[63:0];
    assign _215 = _213[447:64];
    assign _216 = _215[63:0];
    assign _213 = _211[511:64];
    assign _214 = _213[63:0];
    assign _211 = _98[511:0];
    assign _212 = _211[63:0];
    always @* begin
        case (element_offset)
        0: _226 <= _212;
        1: _226 <= _214;
        2: _226 <= _216;
        3: _226 <= _218;
        4: _226 <= _220;
        5: _226 <= _222;
        6: _226 <= _224;
        default: _226 <= _225;
        endcase
    end
    assign _209 = _207[127:64];
    assign _207 = _205[191:64];
    assign _208 = _207[63:0];
    assign _205 = _203[255:64];
    assign _206 = _205[63:0];
    assign _203 = _201[319:64];
    assign _204 = _203[63:0];
    assign _201 = _199[383:64];
    assign _202 = _201[63:0];
    assign _199 = _197[447:64];
    assign _200 = _199[63:0];
    assign _197 = _195[511:64];
    assign _198 = _197[63:0];
    assign _195 = _98[1023:512];
    assign _196 = _195[63:0];
    always @* begin
        case (element_offset)
        0: _210 <= _196;
        1: _210 <= _198;
        2: _210 <= _200;
        3: _210 <= _202;
        4: _210 <= _204;
        5: _210 <= _206;
        6: _210 <= _208;
        default: _210 <= _209;
        endcase
    end
    assign _193 = _191[127:64];
    assign _191 = _189[191:64];
    assign _192 = _191[63:0];
    assign _189 = _187[255:64];
    assign _190 = _189[63:0];
    assign _187 = _185[319:64];
    assign _188 = _187[63:0];
    assign _185 = _183[383:64];
    assign _186 = _185[63:0];
    assign _183 = _181[447:64];
    assign _184 = _183[63:0];
    assign _181 = _179[511:64];
    assign _182 = _181[63:0];
    assign _179 = _98[1535:1024];
    assign _180 = _179[63:0];
    always @* begin
        case (element_offset)
        0: _194 <= _180;
        1: _194 <= _182;
        2: _194 <= _184;
        3: _194 <= _186;
        4: _194 <= _188;
        5: _194 <= _190;
        6: _194 <= _192;
        default: _194 <= _193;
        endcase
    end
    assign _177 = _175[127:64];
    assign _175 = _173[191:64];
    assign _176 = _175[63:0];
    assign _173 = _171[255:64];
    assign _174 = _173[63:0];
    assign _171 = _169[319:64];
    assign _172 = _171[63:0];
    assign _169 = _167[383:64];
    assign _170 = _169[63:0];
    assign _167 = _165[447:64];
    assign _168 = _167[63:0];
    assign _165 = _163[511:64];
    assign _166 = _165[63:0];
    assign _163 = _98[2047:1536];
    assign _164 = _163[63:0];
    always @* begin
        case (element_offset)
        0: _178 <= _164;
        1: _178 <= _166;
        2: _178 <= _168;
        3: _178 <= _170;
        4: _178 <= _172;
        5: _178 <= _174;
        6: _178 <= _176;
        default: _178 <= _177;
        endcase
    end
    assign _161 = _159[127:64];
    assign _159 = _157[191:64];
    assign _160 = _159[63:0];
    assign _157 = _155[255:64];
    assign _158 = _157[63:0];
    assign _155 = _153[319:64];
    assign _156 = _155[63:0];
    assign _153 = _151[383:64];
    assign _154 = _153[63:0];
    assign _151 = _149[447:64];
    assign _152 = _151[63:0];
    assign _149 = _147[511:64];
    assign _150 = _149[63:0];
    assign _147 = _98[2559:2048];
    assign _148 = _147[63:0];
    always @* begin
        case (element_offset)
        0: _162 <= _148;
        1: _162 <= _150;
        2: _162 <= _152;
        3: _162 <= _154;
        4: _162 <= _156;
        5: _162 <= _158;
        6: _162 <= _160;
        default: _162 <= _161;
        endcase
    end
    assign _145 = _143[127:64];
    assign _143 = _141[191:64];
    assign _144 = _143[63:0];
    assign _141 = _139[255:64];
    assign _142 = _141[63:0];
    assign _139 = _137[319:64];
    assign _140 = _139[63:0];
    assign _137 = _135[383:64];
    assign _138 = _137[63:0];
    assign _135 = _133[447:64];
    assign _136 = _135[63:0];
    assign _133 = _131[511:64];
    assign _134 = _133[63:0];
    assign _131 = _98[3071:2560];
    assign _132 = _131[63:0];
    always @* begin
        case (element_offset)
        0: _146 <= _132;
        1: _146 <= _134;
        2: _146 <= _136;
        3: _146 <= _138;
        4: _146 <= _140;
        5: _146 <= _142;
        6: _146 <= _144;
        default: _146 <= _145;
        endcase
    end
    assign _129 = _127[127:64];
    assign _127 = _125[191:64];
    assign _128 = _127[63:0];
    assign _125 = _123[255:64];
    assign _126 = _125[63:0];
    assign _123 = _121[319:64];
    assign _124 = _123[63:0];
    assign _121 = _119[383:64];
    assign _122 = _121[63:0];
    assign _119 = _117[447:64];
    assign _120 = _119[63:0];
    assign _117 = _115[511:64];
    assign _118 = _117[63:0];
    assign _115 = _98[3583:3072];
    assign _116 = _115[63:0];
    always @* begin
        case (element_offset)
        0: _130 <= _116;
        1: _130 <= _118;
        2: _130 <= _120;
        3: _130 <= _122;
        4: _130 <= _124;
        5: _130 <= _126;
        6: _130 <= _128;
        default: _130 <= _129;
        endcase
    end
    assign _113 = _111[127:64];
    assign _111 = _109[191:64];
    assign _112 = _111[63:0];
    assign _109 = _107[255:64];
    assign _110 = _109[63:0];
    assign _107 = _105[319:64];
    assign _108 = _107[63:0];
    assign _105 = _103[383:64];
    assign _106 = _105[63:0];
    assign _103 = _101[447:64];
    assign _104 = _103[63:0];
    assign _101 = _99[511:64];
    assign _102 = _101[63:0];
    assign _11 = in_tdata;
    assign _12 = _11;
    assign _78 = _45 == _42;
    assign _79 = _78 & _22;
    assign _80 = { _79, _79 };
    assign _81 = { _80, _80 };
    assign _82 = { _81, _81 };
    assign _83 = _57 & _82;
    assign _13 = _83;
    assign _84 = _66[0:0];
    assign _85 = { _84, _52 };
    assign _14 = _85;
    assign _89 = _88[0:0];
    assign _93 = { _89, _92 };
    assign _15 = _93;
    transposer_memories
        transposer_memories
        ( .clock(_31), .read_address(_15), .write_address(_14), .write_enable(_13), .write_data(_12), .read_data7(_98[4095:3584]), .read_data6(_98[3583:3072]), .read_data5(_98[3071:2560]), .read_data4(_98[2559:2048]), .read_data3(_98[2047:1536]), .read_data2(_98[1535:1024]), .read_data1(_98[1023:512]), .read_data0(_98[511:0]) );
    assign _99 = _98[4095:3584];
    assign _100 = _99[63:0];
    always @* begin
        case (element_offset)
        0: _114 <= _100;
        1: _114 <= _102;
        2: _114 <= _104;
        3: _114 <= _106;
        4: _114 <= _108;
        5: _114 <= _110;
        6: _114 <= _112;
        default: _114 <= _113;
        endcase
    end
    assign _227 = { _114, _130, _146, _162, _178, _194, _210, _226 };
    assign _16 = _227;
    assign _322 = _308 ? _321 : _315;
    assign _317 = _272 ? _316 : _315;
    assign _318 = _270 ? _317 : _315;
    assign _319 = _34 ? _318 : _315;
    assign _312 = _266 == _267;
    assign _320 = _312 ? _319 : _315;
    assign _306 = wr_pos - _305;
    assign _307 = _88 == _306;
    assign _259 = _66 + _258;
    assign _260 = _58 ? _259 : _66;
    assign _261 = _54 ? _260 : _66;
    assign _262 = _22 ? _261 : _66;
    assign _255 = _71 ? _45 : _42;
    assign _69 = _66 - _68;
    assign _70 = rd_pos == _69;
    assign rd_pos = _88;
    assign _67 = rd_pos == _66;
    assign _71 = _67 | _70;
    assign _240 = _71 ? _239 : _238;
    assign _230 = _57[6:0];
    assign _232 = { _230, _231 };
    assign _234 = _58 ? _233 : _232;
    assign _235 = _54 ? _234 : _57;
    assign _236 = _22 ? _235 : _57;
    assign _229 = _42 == _45;
    assign _237 = _229 ? _236 : _57;
    assign _228 = _42 == _43;
    assign _241 = _228 ? _240 : _237;
    assign _19 = _241;
    always @(posedge _31) begin
        if (_29)
            _57 <= _56;
        else
            _57 <= _19;
    end
    assign _58 = _57[7:7];
    assign _251 = _58 ? _43 : _42;
    assign _244 = _52 + _243;
    assign _246 = _54 ? _245 : _244;
    assign _247 = _22 ? _246 : _52;
    assign _242 = _42 == _45;
    assign _248 = _242 ? _247 : _52;
    assign _20 = _248;
    always @(posedge _31) begin
        if (_29)
            _52 <= _51;
        else
            _52 <= _20;
    end
    assign _54 = _52 == _53;
    assign _252 = _54 ? _251 : _42;
    assign _22 = in_tvalid;
    assign _253 = _22 ? _252 : _42;
    assign _250 = _42 == _45;
    assign _254 = _250 ? _253 : _42;
    assign _249 = _42 == _43;
    assign _256 = _249 ? _255 : _254;
    assign _23 = _256;
    always @(posedge _31) begin
        if (_29)
            _42 <= _40;
        else
            _42 <= _23;
    end
    assign _257 = _42 == _45;
    assign _263 = _257 ? _262 : _66;
    assign _24 = _263;
    always @(posedge _31) begin
        if (_29)
            _66 <= _65;
        else
            _66 <= _24;
    end
    assign wr_pos = _66;
    assign _303 = wr_pos - _302;
    assign _274 = _88 + _273;
    assign _275 = _272 ? _274 : _88;
    assign _276 = _270 ? _275 : _88;
    assign _277 = _34 ? _276 : _88;
    assign _268 = _266 == _267;
    assign _278 = _268 ? _277 : _88;
    assign _26 = _278;
    always @(posedge _31) begin
        if (_29)
            _88 <= _87;
        else
            _88 <= _26;
    end
    assign _304 = _88 == _303;
    assign _308 = _304 | _307;
    assign _309 = _308 ? _267 : _266;
    assign _283 = _92 + _282;
    assign _285 = _272 ? _284 : _283;
    assign _286 = _270 ? _285 : _92;
    assign _287 = _34 ? _286 : _92;
    assign _281 = _266 == _267;
    assign _288 = _281 ? _287 : _92;
    assign _280 = _266 == _279;
    assign _290 = _280 ? _289 : _288;
    assign _27 = _290;
    always @(posedge _31) begin
        if (_29)
            _92 <= _91;
        else
            _92 <= _27;
    end
    assign _272 = _92 == _271;
    assign _298 = _272 ? _279 : _266;
    assign _29 = clear;
    assign _31 = clock;
    assign _293 = element_offset + _292;
    assign _294 = _34 ? _293 : element_offset;
    assign _291 = _266 == _267;
    assign _295 = _291 ? _294 : element_offset;
    assign _32 = _295;
    always @(posedge _31) begin
        if (_29)
            element_offset <= _95;
        else
            element_offset <= _32;
    end
    assign _270 = element_offset == _269;
    assign _299 = _270 ? _298 : _266;
    assign _34 = out_tready;
    assign _300 = _34 ? _299 : _266;
    assign _297 = _266 == _267;
    assign _301 = _297 ? _300 : _266;
    assign _296 = _266 == _279;
    assign _310 = _296 ? _309 : _301;
    assign _35 = _310;
    always @(posedge _31) begin
        if (_29)
            _266 <= _265;
        else
            _266 <= _35;
    end
    assign _311 = _266 == _279;
    assign _323 = _311 ? _322 : _320;
    assign _36 = _323;
    always @(posedge _31) begin
        if (_29)
            _315 <= _314;
        else
            _315 <= _36;
    end
    assign _37 = _315;

    /* aliases */

    /* output assignments */
    assign out_tvalid = _37;
    assign out_tdata = _16;
    assign out_tkeep = _8;
    assign out_tstrb = _6;
    assign out_tlast = _4;
    assign in_tready = _2;

endmodule
module krnl_ntt (
    compute_to_controller_tready,
    controller_to_compute_phase_1_tlast,
    controller_to_compute_phase_1_tstrb,
    controller_to_compute_phase_1_tkeep,
    controller_to_compute_phase_1_tdata,
    controller_to_compute_phase_2_tlast,
    controller_to_compute_phase_2_tstrb,
    controller_to_compute_phase_2_tkeep,
    controller_to_compute_phase_2_tdata,
    controller_to_compute_phase_2_tvalid,
    controller_to_compute_phase_1_tvalid,
    ap_rst_n,
    ap_clk,
    compute_to_controller_tvalid,
    compute_to_controller_tdata,
    compute_to_controller_tkeep,
    compute_to_controller_tstrb,
    compute_to_controller_tlast,
    controller_to_compute_phase_1_tready,
    controller_to_compute_phase_2_tready
);

    input compute_to_controller_tready;
    input controller_to_compute_phase_1_tlast;
    input [63:0] controller_to_compute_phase_1_tstrb;
    input [63:0] controller_to_compute_phase_1_tkeep;
    input [511:0] controller_to_compute_phase_1_tdata;
    input controller_to_compute_phase_2_tlast;
    input [63:0] controller_to_compute_phase_2_tstrb;
    input [63:0] controller_to_compute_phase_2_tkeep;
    input [511:0] controller_to_compute_phase_2_tdata;
    input controller_to_compute_phase_2_tvalid;
    input controller_to_compute_phase_1_tvalid;
    input ap_rst_n;
    input ap_clk;
    output compute_to_controller_tvalid;
    output [511:0] compute_to_controller_tdata;
    output [63:0] compute_to_controller_tkeep;
    output [63:0] compute_to_controller_tstrb;
    output compute_to_controller_tlast;
    output controller_to_compute_phase_1_tready;
    output controller_to_compute_phase_2_tready;

    /* signal declarations */
    wire _41;
    wire _57;
    wire [63:0] _58;
    wire [63:0] _59;
    wire [511:0] _60;
    wire _8;
    wire _10;
    wire _53;
    wire _54;
    wire [63:0] _12;
    wire [63:0] _51;
    wire [63:0] _52;
    wire [63:0] _14;
    wire [63:0] _49;
    wire [63:0] _50;
    wire [511:0] _16;
    wire [511:0] _47;
    wire [511:0] _48;
    wire _61;
    wire _17;
    wire _18;
    wire _20;
    wire [63:0] _22;
    wire [63:0] _24;
    wire [511:0] _26;
    wire [642:0] _40;
    wire _45;
    wire _46;
    wire _43 = 1'b0;
    wire _42 = 1'b0;
    wire _62;
    wire _27;
    reg _4STEP;
    wire _29;
    wire _31;
    wire _64;
    wire _63;
    wire _65;
    wire _32;
    wire _34;
    wire _38;
    wire _36;
    wire [643:0] _56;
    wire _66;

    /* logic */
    assign _41 = _40[642:642];
    assign _57 = _56[641:641];
    assign _58 = _56[640:577];
    assign _59 = _56[576:513];
    assign _60 = _56[512:1];
    assign _8 = compute_to_controller_tready;
    assign _10 = controller_to_compute_phase_1_tlast;
    assign _53 = _40[641:641];
    assign _54 = _31 ? _10 : _53;
    assign _12 = controller_to_compute_phase_1_tstrb;
    assign _51 = _40[640:577];
    assign _52 = _31 ? _12 : _51;
    assign _14 = controller_to_compute_phase_1_tkeep;
    assign _49 = _40[576:513];
    assign _50 = _31 ? _14 : _49;
    assign _16 = controller_to_compute_phase_1_tdata;
    assign _47 = _40[512:1];
    assign _48 = _31 ? _16 : _47;
    assign _61 = _56[642:642];
    assign _17 = _61;
    assign _18 = _17;
    assign _20 = controller_to_compute_phase_2_tlast;
    assign _22 = controller_to_compute_phase_2_tstrb;
    assign _24 = controller_to_compute_phase_2_tkeep;
    assign _26 = controller_to_compute_phase_2_tdata;
    transposer
        transposer
        ( .clock(_36), .clear(_38), .in_tvalid(_29), .in_tdata(_26), .in_tkeep(_24), .in_tstrb(_22), .in_tlast(_20), .out_tready(_18), .in_tready(_40[642:642]), .out_tlast(_40[641:641]), .out_tstrb(_40[640:577]), .out_tkeep(_40[576:513]), .out_tdata(_40[512:1]), .out_tvalid(_40[0:0]) );
    assign _45 = _40[0:0];
    assign _46 = _31 ? _31 : _45;
    assign _62 = ~ _4STEP;
    assign _27 = _62;
    always @(posedge _36) begin
        if (_38)
            _4STEP <= _43;
        else
            if (_32)
                _4STEP <= _27;
    end
    assign _29 = controller_to_compute_phase_2_tvalid;
    assign _31 = controller_to_compute_phase_1_tvalid;
    assign _64 = _31 | _29;
    assign _63 = _56[643:643];
    assign _65 = _63 & _64;
    assign _32 = _65;
    assign _34 = ap_rst_n;
    assign _38 = ~ _34;
    assign _36 = ap_clk;
    kernel
        kernel
        ( .clock(_36), .clear(_38), .start(_32), .first_4step_pass(_4STEP), .data_in_tvalid(_46), .data_in_tdata(_48), .data_in_tkeep(_50), .data_in_tstrb(_52), .data_in_tlast(_54), .data_out_dest_tready(_8), .done_(_56[643:643]), .data_in_dest_tready(_56[642:642]), .data_out_tlast(_56[641:641]), .data_out_tstrb(_56[640:577]), .data_out_tkeep(_56[576:513]), .data_out_tdata(_56[512:1]), .data_out_tvalid(_56[0:0]) );
    assign _66 = _56[0:0];

    /* aliases */

    /* output assignments */
    assign compute_to_controller_tvalid = _66;
    assign compute_to_controller_tdata = _60;
    assign compute_to_controller_tkeep = _59;
    assign compute_to_controller_tstrb = _58;
    assign compute_to_controller_tlast = _57;
    assign controller_to_compute_phase_1_tready = _17;
    assign controller_to_compute_phase_2_tready = _41;

endmodule
