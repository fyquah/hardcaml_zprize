module store_sm (
    start,
    clear,
    clock,
    tready,
    done_,
    tvalid,
    rd_addr,
    rd_en,
    block
);

    input start;
    input clear;
    input clock;
    input tready;
    output done_;
    output tvalid;
    output [11:0] rd_addr;
    output [7:0] rd_en;
    output [2:0] block;

    /* signal declarations */
    wire _56;
    wire _55;
    wire _54;
    wire _52;
    wire _53;
    wire _50;
    wire _51;
    wire _47;
    wire _48;
    wire _49;
    wire _44;
    wire _45;
    wire _46;
    wire _41;
    wire _40;
    wire _42;
    wire [2:0] _24;
    wire _39;
    wire _43;
    wire [7:0] _57;
    wire _33;
    wire _31;
    wire _34;
    wire _29;
    wire _35;
    wire _2;
    wire [1:0] _36;
    wire [3:0] _37;
    wire [7:0] _38;
    wire [7:0] _58;
    wire [14:0] _23;
    wire [11:0] _59;
    wire _63 = 1'b0;
    wire _62 = 1'b0;
    wire _75;
    wire gnd = 1'b0;
    wire _67;
    wire _68;
    wire _61;
    wire _69;
    wire _60;
    wire _76;
    wire _5;
    reg _64;
    wire [1:0] _26 = 2'b00;
    wire [1:0] _25 = 2'b00;
    wire _8;
    wire [1:0] _105;
    wire [3:0] _73 = 4'b1000;
    wire [3:0] _71 = 4'b0000;
    wire [3:0] _70 = 4'b0000;
    wire [3:0] _83 = 4'b0000;
    wire [3:0] _80 = 4'b0001;
    wire [3:0] _81;
    wire _79;
    wire [3:0] _82;
    wire _78;
    wire [3:0] _84;
    wire [3:0] _9;
    reg [3:0] _72;
    wire _74;
    wire [1:0] _103;
    wire [15:0] _65 = 16'b1000000000001000;
    wire vdd = 1'b1;
    wire [15:0] _20 = 16'b0000000000000000;
    wire _11;
    wire [15:0] _19 = 16'b0000000000000000;
    wire _13;
    wire [15:0] _95 = 16'b0000000000000000;
    wire [15:0] _90 = 16'b0000000000000000;
    wire [15:0] _88 = 16'b0000000000000001;
    wire [15:0] _89;
    wire [15:0] _91;
    wire [15:0] _92;
    wire _87;
    wire [15:0] _93;
    wire _86;
    wire [15:0] _94;
    wire _85;
    wire [15:0] _96;
    wire [15:0] _14;
    reg [15:0] _22;
    wire _66;
    wire [1:0] _100;
    wire _16;
    wire [1:0] _101;
    wire [1:0] _30 = 2'b10;
    wire _99;
    wire [1:0] _102;
    wire [1:0] _28 = 2'b01;
    wire _98;
    wire [1:0] _104;
    wire _97;
    wire [1:0] _106;
    wire [1:0] _17;
    reg [1:0] _27;
    wire [1:0] _77 = 2'b00;
    wire _107;

    /* logic */
    assign _56 = _52 & _50;
    assign _55 = _52 & _48;
    assign _54 = _52 & _45;
    assign _52 = ~ _39;
    assign _53 = _52 & _42;
    assign _50 = _47 & _44;
    assign _51 = _39 & _50;
    assign _47 = ~ _40;
    assign _48 = _47 & _41;
    assign _49 = _39 & _48;
    assign _44 = ~ _41;
    assign _45 = _40 & _44;
    assign _46 = _39 & _45;
    assign _41 = _24[0:0];
    assign _40 = _24[1:1];
    assign _42 = _40 & _41;
    assign _24 = _23[2:0];
    assign _39 = _24[2:2];
    assign _43 = _39 & _42;
    assign _57 = { _43, _46, _49, _51, _53, _54, _55, _56 };
    assign _33 = _16 ? vdd : gnd;
    assign _31 = _27 == _30;
    assign _34 = _31 ? _33 : gnd;
    assign _29 = _27 == _28;
    assign _35 = _29 ? vdd : _34;
    assign _2 = _35;
    assign _36 = { _2, _2 };
    assign _37 = { _36, _36 };
    assign _38 = { _37, _37 };
    assign _58 = _38 & _57;
    assign _23 = _22[14:0];
    assign _59 = _23[14:3];
    assign _75 = _74 ? vdd : _64;
    assign _67 = _66 ? gnd : _64;
    assign _68 = _16 ? _67 : _64;
    assign _61 = _27 == _30;
    assign _69 = _61 ? _68 : _64;
    assign _60 = _27 == _28;
    assign _76 = _60 ? _75 : _69;
    assign _5 = _76;
    always @(posedge _13) begin
        if (_11)
            _64 <= _63;
        else
            _64 <= _5;
    end
    assign _8 = start;
    assign _105 = _8 ? _28 : _27;
    assign _81 = _72 + _80;
    assign _79 = _27 == _28;
    assign _82 = _79 ? _81 : _72;
    assign _78 = _27 == _77;
    assign _84 = _78 ? _83 : _82;
    assign _9 = _84;
    always @(posedge _13) begin
        if (_11)
            _72 <= _71;
        else
            _72 <= _9;
    end
    assign _74 = _72 == _73;
    assign _103 = _74 ? _30 : _27;
    assign _11 = clear;
    assign _13 = clock;
    assign _89 = _22 + _88;
    assign _91 = _66 ? _90 : _89;
    assign _92 = _16 ? _91 : _22;
    assign _87 = _27 == _30;
    assign _93 = _87 ? _92 : _22;
    assign _86 = _27 == _28;
    assign _94 = _86 ? _89 : _93;
    assign _85 = _27 == _77;
    assign _96 = _85 ? _95 : _94;
    assign _14 = _96;
    always @(posedge _13) begin
        if (_11)
            _22 <= _20;
        else
            _22 <= _14;
    end
    assign _66 = _22 == _65;
    assign _100 = _66 ? _77 : _27;
    assign _16 = tready;
    assign _101 = _16 ? _100 : _27;
    assign _99 = _27 == _30;
    assign _102 = _99 ? _101 : _27;
    assign _98 = _27 == _28;
    assign _104 = _98 ? _103 : _102;
    assign _97 = _27 == _77;
    assign _106 = _97 ? _105 : _104;
    assign _17 = _106;
    always @(posedge _13) begin
        if (_11)
            _27 <= _26;
        else
            _27 <= _17;
    end
    assign _107 = _77 == _27;

    /* aliases */

    /* output assignments */
    assign done_ = _107;
    assign tvalid = _64;
    assign rd_addr = _59;
    assign rd_en = _58;
    assign block = _24;

endmodule
module controller (
    start,
    clear,
    clock,
    cores_done,
    output_done,
    input_done,
    done_,
    start_input,
    start_output,
    start_cores,
    first_iter,
    flip
);

    input start;
    input clear;
    input clock;
    input cores_done;
    input output_done;
    input input_done;
    output done_;
    output start_input;
    output start_output;
    output start_cores;
    output first_iter;
    output flip;

    /* signal declarations */
    wire _25;
    wire _35 = 1'b1;
    wire _36;
    wire _31;
    wire _37;
    wire _2;
    wire _51;
    wire _48;
    wire _49;
    wire _40;
    wire _50;
    wire _38;
    wire _52;
    wire START_CORES;
    wire _58;
    wire _59;
    wire _56;
    wire _55;
    wire _57;
    wire _53;
    wire _60;
    wire START_OUTPUT;
    wire _70;
    wire _68;
    wire _65;
    wire _66;
    wire gnd = 1'b0;
    wire _64;
    wire _67;
    wire _63;
    wire _69;
    wire _62;
    wire _71;
    wire START_INPUT;
    wire [2:0] _27 = 3'b000;
    wire [2:0] _26 = 3'b000;
    wire _11;
    wire [2:0] _94;
    wire [2:0] _92;
    wire [5:0] _46 = 6'b000000;
    wire [5:0] _44 = 6'b000001;
    wire vdd = 1'b1;
    wire [5:0] _42 = 6'b000000;
    wire _13;
    wire [5:0] _41 = 6'b000000;
    wire _15;
    wire [5:0] _76 = 6'b000001;
    wire [5:0] _77;
    wire [5:0] _74;
    wire _73;
    wire [5:0] _75;
    wire _72;
    wire [5:0] _78;
    wire [5:0] _16;
    reg [5:0] ITERATION;
    wire [5:0] _45;
    wire _47;
    wire [2:0] _89;
    wire [2:0] _90;
    wire [2:0] _87;
    wire _18;
    wire _20;
    wire _22;
    wire _33;
    wire _34;
    wire [2:0] _85;
    wire [2:0] _83 = 3'b100;
    wire _84;
    wire [2:0] _86;
    wire [2:0] _54 = 3'b011;
    wire _82;
    wire [2:0] _88;
    wire [2:0] _39 = 3'b010;
    wire _81;
    wire [2:0] _91;
    wire [2:0] _30 = 3'b001;
    wire _80;
    wire [2:0] _93;
    wire _79;
    wire [2:0] _95;
    wire [2:0] _23;
    reg [2:0] STATE;
    wire [2:0] _61 = 3'b000;
    wire _96;

    /* logic */
    assign _25 = START_CORES | START_OUTPUT;
    assign _36 = _34 ? _35 : gnd;
    assign _31 = STATE == _30;
    assign _37 = _31 ? _36 : gnd;
    assign _2 = _37;
    assign _51 = _34 ? vdd : gnd;
    assign _48 = _47 ? vdd : vdd;
    assign _49 = _34 ? _48 : gnd;
    assign _40 = STATE == _39;
    assign _50 = _40 ? _49 : gnd;
    assign _38 = STATE == _30;
    assign _52 = _38 ? _51 : _50;
    assign START_CORES = _52;
    assign _58 = _47 ? vdd : vdd;
    assign _59 = _34 ? _58 : gnd;
    assign _56 = _34 ? vdd : gnd;
    assign _55 = STATE == _54;
    assign _57 = _55 ? _56 : gnd;
    assign _53 = STATE == _39;
    assign _60 = _53 ? _59 : _57;
    assign START_OUTPUT = _60;
    assign _70 = _11 ? vdd : gnd;
    assign _68 = _34 ? vdd : gnd;
    assign _65 = _47 ? gnd : vdd;
    assign _66 = _34 ? _65 : gnd;
    assign _64 = STATE == _39;
    assign _67 = _64 ? _66 : gnd;
    assign _63 = STATE == _30;
    assign _69 = _63 ? _68 : _67;
    assign _62 = STATE == _61;
    assign _71 = _62 ? _70 : _69;
    assign START_INPUT = _71;
    assign _11 = start;
    assign _94 = _11 ? _30 : STATE;
    assign _92 = _34 ? _39 : STATE;
    assign _13 = clear;
    assign _15 = clock;
    assign _77 = _34 ? _76 : ITERATION;
    assign _74 = _34 ? _45 : ITERATION;
    assign _73 = STATE == _39;
    assign _75 = _73 ? _74 : ITERATION;
    assign _72 = STATE == _30;
    assign _78 = _72 ? _77 : _75;
    assign _16 = _78;
    always @(posedge _15) begin
        if (_13)
            ITERATION <= _42;
        else
            ITERATION <= _16;
    end
    assign _45 = ITERATION + _44;
    assign _47 = _45 == _46;
    assign _89 = _47 ? _54 : STATE;
    assign _90 = _34 ? _89 : STATE;
    assign _87 = _34 ? _83 : STATE;
    assign _18 = cores_done;
    assign _20 = output_done;
    assign _22 = input_done;
    assign _33 = _22 & _20;
    assign _34 = _33 & _18;
    assign _85 = _34 ? _61 : STATE;
    assign _84 = STATE == _83;
    assign _86 = _84 ? _85 : STATE;
    assign _82 = STATE == _54;
    assign _88 = _82 ? _87 : _86;
    assign _81 = STATE == _39;
    assign _91 = _81 ? _90 : _88;
    assign _80 = STATE == _30;
    assign _93 = _80 ? _92 : _91;
    assign _79 = STATE == _61;
    assign _95 = _79 ? _94 : _93;
    assign _23 = _95;
    always @(posedge _15) begin
        if (_13)
            STATE <= _27;
        else
            STATE <= _23;
    end
    assign _96 = _61 == STATE;

    /* aliases */

    /* output assignments */
    assign done_ = _96;
    assign start_input = START_INPUT;
    assign start_output = START_OUTPUT;
    assign start_cores = START_CORES;
    assign first_iter = _2;
    assign flip = _25;

endmodule
module load_sm (
    first_4step_pass,
    start,
    tvalid,
    clear,
    clock,
    done_,
    tready,
    wr_addr,
    wr_en
);

    input first_4step_pass;
    input start;
    input tvalid;
    input clear;
    input clock;
    output done_;
    output tready;
    output [11:0] wr_addr;
    output [7:0] wr_en;

    /* signal declarations */
    wire _51;
    wire _50;
    wire _49;
    wire _47;
    wire _48;
    wire _45;
    wire _46;
    wire _42;
    wire _43;
    wire _44;
    wire _39;
    wire _40;
    wire _41;
    wire _36;
    wire _35;
    wire _37;
    wire [2:0] _32;
    wire [2:0] _31;
    wire [2:0] _33;
    wire _34;
    wire _38;
    wire [7:0] _52;
    wire _24;
    wire [1:0] _25;
    wire [3:0] _26;
    wire [7:0] _27;
    wire [7:0] _53;
    wire [11:0] _55;
    wire [11:0] _54;
    wire _3;
    wire [11:0] _56;
    wire _23;
    wire [1:0] _20 = 2'b00;
    wire [1:0] _19 = 2'b00;
    wire _7;
    wire [1:0] _89;
    wire [14:0] _84 = 15'b000000000000000;
    wire [14:0] _60 = 15'b000000000000001;
    wire [14:0] _29 = 15'b000000000000000;
    wire [14:0] _28 = 15'b000000000000000;
    wire [14:0] _64 = 15'b000000000000000;
    wire [14:0] _62;
    wire _59;
    wire [14:0] _63;
    wire _58;
    wire [14:0] _65;
    wire [14:0] _8;
    reg [14:0] _30;
    wire [14:0] _61;
    wire _85;
    wire [1:0] _86;
    wire _10;
    wire [1:0] _87;
    wire _80 = 1'b1;
    wire vdd = 1'b1;
    wire _70 = 1'b0;
    wire _12;
    wire _69 = 1'b0;
    wire _14;
    wire _75 = 1'b0;
    wire _72 = 1'b1;
    wire _73;
    wire _68;
    wire _74;
    wire _66;
    wire _76;
    wire _15;
    reg _71;
    wire _81;
    wire [1:0] _82;
    wire [1:0] _67 = 2'b10;
    wire _79;
    wire [1:0] _83;
    wire [1:0] _18 = 2'b01;
    wire _78;
    wire [1:0] _88;
    wire _77;
    wire [1:0] _90;
    wire [1:0] _16;
    reg [1:0] _22;
    wire [1:0] _57 = 2'b00;
    wire _91;

    /* logic */
    assign _51 = _47 & _45;
    assign _50 = _47 & _43;
    assign _49 = _47 & _40;
    assign _47 = ~ _34;
    assign _48 = _47 & _37;
    assign _45 = _42 & _39;
    assign _46 = _34 & _45;
    assign _42 = ~ _35;
    assign _43 = _42 & _36;
    assign _44 = _34 & _43;
    assign _39 = ~ _36;
    assign _40 = _35 & _39;
    assign _41 = _34 & _40;
    assign _36 = _33[0:0];
    assign _35 = _33[1:1];
    assign _37 = _35 & _36;
    assign _32 = _30[2:0];
    assign _31 = _30[14:12];
    assign _33 = _3 ? _32 : _31;
    assign _34 = _33[2:2];
    assign _38 = _34 & _37;
    assign _52 = { _38, _41, _44, _46, _48, _49, _50, _51 };
    assign _24 = _23 & _10;
    assign _25 = { _24, _24 };
    assign _26 = { _25, _25 };
    assign _27 = { _26, _26 };
    assign _53 = _27 & _52;
    assign _55 = _30[14:3];
    assign _54 = _30[11:0];
    assign _3 = first_4step_pass;
    assign _56 = _3 ? _55 : _54;
    assign _23 = _18 == _22;
    assign _7 = start;
    assign _89 = _7 ? _18 : _22;
    assign _62 = _10 ? _61 : _30;
    assign _59 = _22 == _18;
    assign _63 = _59 ? _62 : _30;
    assign _58 = _22 == _57;
    assign _65 = _58 ? _64 : _63;
    assign _8 = _65;
    always @(posedge _14) begin
        if (_12)
            _30 <= _29;
        else
            _30 <= _8;
    end
    assign _61 = _30 + _60;
    assign _85 = _61 == _84;
    assign _86 = _85 ? _67 : _22;
    assign _10 = tvalid;
    assign _87 = _10 ? _86 : _22;
    assign _12 = clear;
    assign _14 = clock;
    assign _73 = _71 + _72;
    assign _68 = _22 == _67;
    assign _74 = _68 ? _73 : _71;
    assign _66 = _22 == _57;
    assign _76 = _66 ? _75 : _74;
    assign _15 = _76;
    always @(posedge _14) begin
        if (_12)
            _71 <= _70;
        else
            _71 <= _15;
    end
    assign _81 = _71 == _80;
    assign _82 = _81 ? _57 : _22;
    assign _79 = _22 == _67;
    assign _83 = _79 ? _82 : _22;
    assign _78 = _22 == _18;
    assign _88 = _78 ? _87 : _83;
    assign _77 = _22 == _57;
    assign _90 = _77 ? _89 : _88;
    assign _16 = _90;
    always @(posedge _14) begin
        if (_12)
            _22 <= _20;
        else
            _22 <= _16;
    end
    assign _91 = _57 == _22;

    /* aliases */

    /* output assignments */
    assign done_ = _91;
    assign tready = _23;
    assign wr_addr = _56;
    assign wr_en = _53;

endmodule
module ctrl (
    first_4step_pass,
    start,
    clear,
    clock,
    first_iter,
    done_,
    i,
    j,
    k,
    m,
    addr1,
    addr2,
    omegas0,
    omegas1,
    omegas2,
    omegas3,
    omegas4,
    omegas5,
    omegas6,
    start_twiddles,
    first_stage,
    last_stage,
    twiddle_stage,
    valid,
    index,
    read_write_enable,
    flip
);

    input first_4step_pass;
    input start;
    input clear;
    input clock;
    input first_iter;
    output done_;
    output [3:0] i;
    output [11:0] j;
    output [11:0] k;
    output [11:0] m;
    output [11:0] addr1;
    output [11:0] addr2;
    output [63:0] omegas0;
    output [63:0] omegas1;
    output [63:0] omegas2;
    output [63:0] omegas3;
    output [63:0] omegas4;
    output [63:0] omegas5;
    output [63:0] omegas6;
    output start_twiddles;
    output first_stage;
    output last_stage;
    output twiddle_stage;
    output valid;
    output [3:0] index;
    output read_write_enable;
    output flip;

    /* signal declarations */
    wire _59;
    wire _52;
    wire _60;
    wire _1;
    wire _64;
    wire _65;
    wire _62;
    wire _66;
    wire _3;
    wire _73 = 1'b0;
    wire _72 = 1'b0;
    wire _92 = 1'b0;
    wire _93;
    wire _89 = 1'b1;
    wire _90;
    wire _81 = 1'b0;
    wire _79 = 1'b0;
    wire [3:0] _77 = 4'b0110;
    wire _78;
    wire _80;
    wire _82;
    wire _71;
    wire _83;
    wire _69;
    wire _91;
    wire _68;
    wire _94;
    wire _6;
    reg _74;
    wire _100 = 1'b0;
    wire _99 = 1'b0;
    wire _120 = 1'b0;
    wire _121;
    wire _115 = 1'b1;
    wire _116;
    wire _117;
    wire _118;
    wire _105 = 1'b0;
    wire _106;
    wire _102 = 1'b0;
    wire _103;
    wire _98;
    wire _104;
    wire _97;
    wire _107;
    wire _96;
    wire _119;
    wire _95;
    wire _122;
    wire _8;
    reg _101;
    wire _127 = 1'b0;
    wire _126 = 1'b0;
    wire _141 = 1'b0;
    wire _142;
    wire _136 = 1'b1;
    wire _135 = 1'b0;
    wire _137;
    wire _133;
    wire [3:0] _131 = 4'b1011;
    wire _132;
    wire _134;
    wire _138;
    wire _139;
    wire gnd = 1'b0;
    wire _129;
    wire _125;
    wire _130;
    wire _124;
    wire _140;
    wire _123;
    wire _143;
    wire _10;
    reg _128;
    wire _147 = 1'b0;
    wire _146 = 1'b0;
    wire _152 = 1'b1;
    wire _153;
    wire _149 = 1'b0;
    wire _150;
    wire _145;
    wire _151;
    wire _144;
    wire _154;
    wire _12;
    reg _148;
    wire _188 = 1'b0;
    wire _187 = 1'b0;
    wire _184 = 1'b1;
    wire _185;
    wire _180 = 1'b1;
    wire _181;
    wire _182;
    wire _159 = 1'b1;
    wire _160;
    wire _158 = 1'b0;
    wire _157;
    wire _161;
    wire _156;
    wire _183;
    wire _155;
    wire _186;
    wire _14;
    reg _189;
    wire [63:0] _201 = 64'b1110000010010110111101100111110101000010010111011100100100000111;
    wire [63:0] _200 = 64'b1110111110011011001000010110000110000111101001101001011101000111;
    wire [63:0] _199 = 64'b0101010011010111101011100001010011111111011110000011001100001001;
    wire [63:0] _198 = 64'b1001010110000011011011011110011100001111001100011100101111111010;
    wire [63:0] _197 = 64'b0011101110101011111110001010011100001011100100000001011011010111;
    wire [63:0] _196 = 64'b1111111111111111111111111111110111111111111111110000000000000010;
    wire [63:0] _195 = 64'b0000000000000001111111111111111111111111111111100000000000000000;
    wire [63:0] _194 = 64'b1111111111111111111111111111101100000000000000000000000000000101;
    wire [63:0] _193 = 64'b1111111111111111111111111110111100000000000000000000000000000001;
    wire [63:0] _192 = 64'b0000000000000000000000001111111111111111111111111111111100000000;
    wire [63:0] _191 = 64'b1111111111111110111111111111111100000000000000000000000000000001;
    wire [63:0] _190 = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    reg [63:0] _202;
    wire [63:0] _214 = 64'b0110111000001001111101011111101101111110101000111110001001000001;
    wire [63:0] _213 = 64'b0110000010000100111001101000010001011010100100010010111101001101;
    wire [63:0] _212 = 64'b1011101000100101111010110101110011010001100101110000101011101011;
    wire [63:0] _211 = 64'b0000001111101000110111111101001001001110100011100111100000011111;
    wire [63:0] _210 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _209 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _208 = 64'b0000000000000000000001000000000000000000000000000000000000000000;
    wire [63:0] _207 = 64'b0000000000001111111111111111111111111111111100000000000000000000;
    wire [63:0] _206 = 64'b1111111111111111111111101111111100000000000000000000000100000001;
    wire [63:0] _205 = 64'b1111111111111110111111111111111100000000000000000000000000000001;
    wire [63:0] _204 = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [63:0] _203 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    reg [63:0] _215;
    wire [63:0] _227 = 64'b1001100001001110110001010001100101001101000000000101011100110101;
    wire [63:0] _226 = 64'b0111101001011001000101011001010111100110011111000010011111101000;
    wire [63:0] _225 = 64'b0011110110100000010111111110111001110000110001001111001010111010;
    wire [63:0] _224 = 64'b1100100001000011111100010110001010010100011000001011010101010001;
    wire [63:0] _223 = 64'b1100001011011110110100010111001001000011011101011110000100101110;
    wire [63:0] _222 = 64'b0000000000000000000000011111111111111101111111111111111000000000;
    wire [63:0] _221 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
    wire [63:0] _220 = 64'b0000000000000000000000000000000000000000000000000000000001000000;
    wire [63:0] _219 = 64'b0000000000000000000000000000000000000000000000000001000000000000;
    wire [63:0] _218 = 64'b0000000000000000000000000000000000000001000000000000000000000000;
    wire [63:0] _217 = 64'b0000000000000001000000000000000000000000000000000000000000000000;
    wire [63:0] _216 = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    reg [63:0] _228;
    wire [63:0] _240 = 64'b1001110110001111001010101101011110001011111111101101100101110010;
    wire [63:0] _239 = 64'b0001100100000101110100000010101001011100010000010001111101001110;
    wire [63:0] _238 = 64'b1011111101111001000101000011110011100110000011001010100101100110;
    wire [63:0] _237 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    wire [63:0] _236 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _234 = 64'b1110111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _233 = 64'b1111111111111111111111111111111011111111000000000000000000000001;
    wire [63:0] _232 = 64'b0000000000000001000000000000000000000000000000000000000000000000;
    wire [63:0] _231 = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [63:0] _230 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _229 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    reg [63:0] _241;
    wire [63:0] _253 = 64'b1001010001011000110101001011010000001101001101000000011100011110;
    wire [63:0] _252 = 64'b0110111000001001111101011111101101111110101000111110001001000001;
    wire [63:0] _251 = 64'b0110000010000100111001101000010001011010100100010010111101001101;
    wire [63:0] _250 = 64'b1011101000100101111010110101110011010001100101110000101011101011;
    wire [63:0] _249 = 64'b0000001111101000110111111101001001001110100011100111100000011111;
    wire [63:0] _248 = 64'b0000000000000100000000000000001111111111111111000000000000000000;
    wire [63:0] _247 = 64'b1111111111111111111111111111111011111111111000000000000000000001;
    wire [63:0] _246 = 64'b0000000000000000000001000000000000000000000000000000000000000000;
    wire [63:0] _245 = 64'b0000000000001111111111111111111111111111111100000000000000000000;
    wire [63:0] _244 = 64'b1111111111111111111111101111111100000000000000000000000100000001;
    wire [63:0] _243 = 64'b1111111111111110111111111111111100000000000000000000000000000001;
    wire [63:0] _242 = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    reg [63:0] _254;
    wire [63:0] _266 = 64'b0000011001010011101101001000000000011101101000011100100011001111;
    wire [63:0] _265 = 64'b1001110110001111001010101101011110001011111111101101100101110010;
    wire [63:0] _264 = 64'b0001100100000101110100000010101001011100010000010001111101001110;
    wire [63:0] _263 = 64'b1011111101111001000101000011110011100110000011001010100101100110;
    wire [63:0] _262 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    wire [63:0] _261 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _260 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _259 = 64'b1110111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _258 = 64'b1111111111111111111111111111111011111111000000000000000000000001;
    wire [63:0] _257 = 64'b0000000000000001000000000000000000000000000000000000000000000000;
    wire [63:0] _256 = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    wire [63:0] _255 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    reg [63:0] _267;
    wire [63:0] _279 = 64'b1111001011000011010100011001100110010101100111011111110010110110;
    wire [63:0] _278 = 64'b0000011001010011101101001000000000011101101000011100100011001111;
    wire [63:0] _277 = 64'b1001110110001111001010101101011110001011111111101101100101110010;
    wire [63:0] _276 = 64'b0001100100000101110100000010101001011100010000010001111101001110;
    wire [63:0] _275 = 64'b1011111101111001000101000011110011100110000011001010100101100110;
    wire [63:0] _274 = 64'b1111100000000000000001111111111100001000000000000000000000000001;
    wire [63:0] _273 = 64'b0000000000000000000000001000000000000000000000000000000000000000;
    wire [63:0] _272 = 64'b0000000000000000001111111111111111111111111111111100000000000000;
    wire [63:0] _271 = 64'b1110111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _270 = 64'b1111111111111111111111111111111011111111000000000000000000000001;
    wire [63:0] _269 = 64'b0000000000000001000000000000000000000000000000000000000000000000;
    wire [63:0] _268 = 64'b1111111111111111111111111111111100000000000000000000000000000000;
    reg [63:0] _280;
    wire [11:0] _285 = 12'b000000000000;
    wire [11:0] _284 = 12'b000000000000;
    wire [11:0] _294 = 12'b000000000000;
    wire [11:0] _295;
    wire [11:0] _291;
    wire [11:0] _289 = 12'b000000000001;
    wire [11:0] _290;
    wire [11:0] _292;
    wire [11:0] _287;
    wire _283;
    wire [11:0] _288;
    wire _282;
    wire [11:0] _293;
    wire _281;
    wire [11:0] _296;
    wire [11:0] _24;
    reg [11:0] _286;
    wire _386 = 1'b0;
    wire _396 = 1'b0;
    wire _397;
    wire _391 = 1'b1;
    wire _392;
    wire _393;
    wire _394;
    wire _388 = 1'b1;
    wire _389;
    wire _385;
    wire _390;
    wire _384;
    wire _395;
    wire [2:0] _48 = 3'b000;
    wire [2:0] _47 = 3'b000;
    wire [2:0] _381;
    wire [2:0] _378;
    wire [2:0] _379;
    wire [2:0] _374;
    wire [2:0] _375;
    wire [2:0] _376;
    wire [11:0] _87 = 12'b111111111111;
    wire [11:0] _85 = 12'b000000000000;
    wire [11:0] _84 = 12'b000000000000;
    wire [11:0] _354 = 12'b000000000001;
    wire [11:0] _355;
    wire [11:0] _350;
    wire [11:0] _351;
    wire [11:0] _352;
    wire [11:0] _345 = 12'b000000000000;
    wire _31;
    wire [11:0] _346;
    wire [11:0] _172 = 12'b000000000000;
    wire [11:0] _171 = 12'b000000000000;
    wire [11:0] _325 = 12'b000000000000;
    wire [11:0] _326;
    wire [11:0] _322;
    wire [11:0] _168 = 12'b000000000000;
    wire [11:0] _167 = 12'b000000000000;
    wire [11:0] _301 = 12'b000000000001;
    wire [11:0] _302;
    wire _175 = 1'b0;
    wire [10:0] _174;
    wire [11:0] _176;
    wire [11:0] _299;
    wire _298;
    wire [11:0] _300;
    wire _297;
    wire [11:0] _303;
    wire [11:0] _32;
    reg [11:0] m_0;
    wire [11:0] _165 = 12'b000000000001;
    wire [11:0] _163 = 12'b000000000000;
    wire [11:0] _162 = 12'b000000000000;
    wire [11:0] _314 = 12'b000000000000;
    wire [11:0] _315;
    wire [11:0] _310 = 12'b000000000000;
    wire [11:0] _178 = 12'b000000000000;
    wire _179;
    wire [11:0] _311;
    wire [11:0] _312;
    wire [11:0] _307 = 12'b000000000000;
    wire [11:0] _308;
    wire _306;
    wire [11:0] _309;
    wire _305;
    wire [11:0] _313;
    wire _304;
    wire [11:0] _316;
    wire [11:0] _33;
    reg [11:0] j_0;
    wire [11:0] _166;
    wire _170;
    wire [11:0] _323;
    wire [11:0] _320;
    wire _319;
    wire [11:0] _321;
    wire _318;
    wire [11:0] _324;
    wire _317;
    wire [11:0] _327;
    wire [11:0] _34;
    reg [11:0] k_0;
    wire [11:0] _177;
    wire [11:0] _344;
    wire [3:0] _113 = 4'b1100;
    wire [3:0] _111 = 4'b0001;
    wire [3:0] _109 = 4'b0000;
    wire [3:0] _108 = 4'b0000;
    wire [3:0] _332 = 4'b0000;
    wire _36;
    wire [3:0] _333;
    wire [3:0] _330;
    wire _329;
    wire [3:0] _331;
    wire _328;
    wire [3:0] _334;
    wire [3:0] _37;
    reg [3:0] i_0;
    wire [3:0] _112;
    wire _114;
    wire [11:0] _347;
    wire [11:0] _348;
    wire [11:0] _341 = 12'b000000000000;
    wire [11:0] _339 = 12'b000000000001;
    wire [11:0] _340;
    wire [11:0] _342;
    wire _338;
    wire [11:0] _343;
    wire _337;
    wire [11:0] _349;
    wire _336;
    wire [11:0] _353;
    wire _335;
    wire [11:0] _356;
    wire [11:0] _38;
    reg [11:0] _86;
    wire _88;
    wire [2:0] _372;
    wire [3:0] _75 = 4'b1000;
    wire vdd = 1'b1;
    wire [3:0] _55 = 4'b0000;
    wire _40;
    wire [3:0] _54 = 4'b0000;
    wire _42;
    wire [3:0] _362 = 4'b0000;
    wire [3:0] _57 = 4'b1000;
    wire _58;
    wire [3:0] _363;
    wire [3:0] _359 = 4'b0001;
    wire [3:0] _360;
    wire _358;
    wire [3:0] _361;
    wire _357;
    wire [3:0] _364;
    wire [3:0] _43;
    reg [3:0] _56;
    wire _76;
    wire [2:0] _370;
    wire [2:0] _70 = 3'b100;
    wire _369;
    wire [2:0] _371;
    wire [2:0] _63 = 3'b011;
    wire _368;
    wire [2:0] _373;
    wire [2:0] _51 = 3'b010;
    wire _367;
    wire [2:0] _377;
    wire [2:0] _61 = 3'b001;
    wire _366;
    wire [2:0] _380;
    wire [2:0] _67 = 3'b000;
    wire _365;
    wire [2:0] _382;
    wire [2:0] _44;
    reg [2:0] STATE;
    wire _383;
    wire _398;
    wire _45;
    reg _387;

    /* logic */
    assign _59 = _58 ? vdd : gnd;
    assign _52 = STATE == _51;
    assign _60 = _52 ? _59 : gnd;
    assign _1 = _60;
    assign _64 = STATE == _63;
    assign _65 = _64 ? vdd : gnd;
    assign _62 = STATE == _61;
    assign _66 = _62 ? vdd : _65;
    assign _3 = _66;
    assign _93 = _36 ? _92 : _74;
    assign _90 = _88 ? _89 : _74;
    assign _78 = _56 == _77;
    assign _80 = _78 ? _79 : _74;
    assign _82 = _76 ? _81 : _80;
    assign _71 = STATE == _70;
    assign _83 = _71 ? _82 : _74;
    assign _69 = STATE == _63;
    assign _91 = _69 ? _90 : _83;
    assign _68 = STATE == _67;
    assign _94 = _68 ? _93 : _91;
    assign _6 = _94;
    always @(posedge _42) begin
        if (_40)
            _74 <= _73;
        else
            _74 <= _6;
    end
    assign _121 = _36 ? _120 : _101;
    assign _116 = _31 ? _115 : _101;
    assign _117 = _114 ? _116 : _101;
    assign _118 = _58 ? _117 : _101;
    assign _106 = _88 ? _105 : _101;
    assign _103 = _76 ? _102 : _101;
    assign _98 = STATE == _70;
    assign _104 = _98 ? _103 : _101;
    assign _97 = STATE == _63;
    assign _107 = _97 ? _106 : _104;
    assign _96 = STATE == _51;
    assign _119 = _96 ? _118 : _107;
    assign _95 = STATE == _67;
    assign _122 = _95 ? _121 : _119;
    assign _8 = _122;
    always @(posedge _42) begin
        if (_40)
            _101 <= _100;
        else
            _101 <= _8;
    end
    assign _142 = _36 ? _141 : _128;
    assign _137 = _31 ? _136 : _135;
    assign _133 = ~ _31;
    assign _132 = _112 == _131;
    assign _134 = _132 ? _133 : _128;
    assign _138 = _114 ? _137 : _134;
    assign _139 = _58 ? _138 : _128;
    assign _129 = _76 ? gnd : _128;
    assign _125 = STATE == _70;
    assign _130 = _125 ? _129 : _128;
    assign _124 = STATE == _51;
    assign _140 = _124 ? _139 : _130;
    assign _123 = STATE == _67;
    assign _143 = _123 ? _142 : _140;
    assign _10 = _143;
    always @(posedge _42) begin
        if (_40)
            _128 <= _127;
        else
            _128 <= _10;
    end
    assign _153 = _36 ? _152 : _148;
    assign _150 = _58 ? _149 : _148;
    assign _145 = STATE == _51;
    assign _151 = _145 ? _150 : _148;
    assign _144 = STATE == _67;
    assign _154 = _144 ? _153 : _151;
    assign _12 = _154;
    always @(posedge _42) begin
        if (_40)
            _148 <= _147;
        else
            _148 <= _12;
    end
    assign _185 = _36 ? _184 : _158;
    assign _181 = _179 ? _158 : _180;
    assign _182 = _170 ? _181 : _158;
    assign _160 = _58 ? _159 : _158;
    assign _157 = STATE == _51;
    assign _161 = _157 ? _160 : _158;
    assign _156 = STATE == _61;
    assign _183 = _156 ? _182 : _161;
    assign _155 = STATE == _67;
    assign _186 = _155 ? _185 : _183;
    assign _14 = _186;
    always @(posedge _42) begin
        if (_40)
            _189 <= _188;
        else
            _189 <= _14;
    end
    always @* begin
        case (i_0)
        0: _202 <= _190;
        1: _202 <= _191;
        2: _202 <= _192;
        3: _202 <= _193;
        4: _202 <= _194;
        5: _202 <= _195;
        6: _202 <= _196;
        7: _202 <= _197;
        8: _202 <= _198;
        9: _202 <= _199;
        10: _202 <= _200;
        default: _202 <= _201;
        endcase
    end
    always @* begin
        case (i_0)
        0: _215 <= _203;
        1: _215 <= _204;
        2: _215 <= _205;
        3: _215 <= _206;
        4: _215 <= _207;
        5: _215 <= _208;
        6: _215 <= _209;
        7: _215 <= _210;
        8: _215 <= _211;
        9: _215 <= _212;
        10: _215 <= _213;
        default: _215 <= _214;
        endcase
    end
    always @* begin
        case (i_0)
        0: _228 <= _216;
        1: _228 <= _217;
        2: _228 <= _218;
        3: _228 <= _219;
        4: _228 <= _220;
        5: _228 <= _221;
        6: _228 <= _222;
        7: _228 <= _223;
        8: _228 <= _224;
        9: _228 <= _225;
        10: _228 <= _226;
        default: _228 <= _227;
        endcase
    end
    always @* begin
        case (i_0)
        0: _241 <= _229;
        1: _241 <= _230;
        2: _241 <= _231;
        3: _241 <= _232;
        4: _241 <= _233;
        5: _241 <= _234;
        6: _241 <= _235;
        7: _241 <= _236;
        8: _241 <= _237;
        9: _241 <= _238;
        10: _241 <= _239;
        default: _241 <= _240;
        endcase
    end
    always @* begin
        case (i_0)
        0: _254 <= _242;
        1: _254 <= _243;
        2: _254 <= _244;
        3: _254 <= _245;
        4: _254 <= _246;
        5: _254 <= _247;
        6: _254 <= _248;
        7: _254 <= _249;
        8: _254 <= _250;
        9: _254 <= _251;
        10: _254 <= _252;
        default: _254 <= _253;
        endcase
    end
    always @* begin
        case (i_0)
        0: _267 <= _255;
        1: _267 <= _256;
        2: _267 <= _257;
        3: _267 <= _258;
        4: _267 <= _259;
        5: _267 <= _260;
        6: _267 <= _261;
        7: _267 <= _262;
        8: _267 <= _263;
        9: _267 <= _264;
        10: _267 <= _265;
        default: _267 <= _266;
        endcase
    end
    always @* begin
        case (i_0)
        0: _280 <= _268;
        1: _280 <= _269;
        2: _280 <= _270;
        3: _280 <= _271;
        4: _280 <= _272;
        5: _280 <= _273;
        6: _280 <= _274;
        7: _280 <= _275;
        8: _280 <= _276;
        9: _280 <= _277;
        10: _280 <= _278;
        default: _280 <= _279;
        endcase
    end
    assign _295 = _36 ? _294 : _286;
    assign _291 = _179 ? _290 : _177;
    assign _290 = _286 + _289;
    assign _292 = _170 ? _291 : _290;
    assign _287 = _58 ? _177 : _286;
    assign _283 = STATE == _51;
    assign _288 = _283 ? _287 : _286;
    assign _282 = STATE == _61;
    assign _293 = _282 ? _292 : _288;
    assign _281 = STATE == _67;
    assign _296 = _281 ? _295 : _293;
    assign _24 = _296;
    always @(posedge _42) begin
        if (_40)
            _286 <= _285;
        else
            _286 <= _24;
    end
    assign _397 = _36 ? _396 : _387;
    assign _392 = _31 ? _387 : _391;
    assign _393 = _114 ? _392 : _387;
    assign _394 = _58 ? _393 : _387;
    assign _389 = _76 ? _388 : _387;
    assign _385 = STATE == _70;
    assign _390 = _385 ? _389 : _387;
    assign _384 = STATE == _51;
    assign _395 = _384 ? _394 : _390;
    assign _381 = _36 ? _61 : STATE;
    assign _378 = _179 ? _51 : STATE;
    assign _379 = _170 ? _378 : STATE;
    assign _374 = _31 ? _63 : _67;
    assign _375 = _114 ? _374 : _61;
    assign _376 = _58 ? _375 : STATE;
    assign _355 = _36 ? _354 : _86;
    assign _350 = _177 + m_0;
    assign _351 = _179 ? _340 : _350;
    assign _352 = _170 ? _351 : _340;
    assign _31 = first_4step_pass;
    assign _346 = _31 ? _345 : _344;
    assign _326 = _36 ? _325 : k_0;
    assign _322 = _179 ? k_0 : _177;
    assign _302 = _36 ? _301 : m_0;
    assign _174 = m_0[10:0];
    assign _176 = { _174, _175 };
    assign _299 = _58 ? _176 : m_0;
    assign _298 = STATE == _51;
    assign _300 = _298 ? _299 : m_0;
    assign _297 = STATE == _67;
    assign _303 = _297 ? _302 : _300;
    assign _32 = _303;
    always @(posedge _42) begin
        if (_40)
            m_0 <= _168;
        else
            m_0 <= _32;
    end
    assign _315 = _36 ? _314 : j_0;
    assign _179 = _177 == _178;
    assign _311 = _179 ? _166 : _310;
    assign _312 = _170 ? _311 : _166;
    assign _308 = _58 ? _307 : j_0;
    assign _306 = STATE == _51;
    assign _309 = _306 ? _308 : j_0;
    assign _305 = STATE == _61;
    assign _313 = _305 ? _312 : _309;
    assign _304 = STATE == _67;
    assign _316 = _304 ? _315 : _313;
    assign _33 = _316;
    always @(posedge _42) begin
        if (_40)
            j_0 <= _163;
        else
            j_0 <= _33;
    end
    assign _166 = j_0 + _165;
    assign _170 = _166 == m_0;
    assign _323 = _170 ? _322 : k_0;
    assign _320 = _58 ? _177 : k_0;
    assign _319 = STATE == _51;
    assign _321 = _319 ? _320 : k_0;
    assign _318 = STATE == _61;
    assign _324 = _318 ? _323 : _321;
    assign _317 = STATE == _67;
    assign _327 = _317 ? _326 : _324;
    assign _34 = _327;
    always @(posedge _42) begin
        if (_40)
            k_0 <= _172;
        else
            k_0 <= _34;
    end
    assign _177 = k_0 + _176;
    assign _344 = _177 + _176;
    assign _36 = start;
    assign _333 = _36 ? _332 : i_0;
    assign _330 = _58 ? _112 : i_0;
    assign _329 = STATE == _51;
    assign _331 = _329 ? _330 : i_0;
    assign _328 = STATE == _67;
    assign _334 = _328 ? _333 : _331;
    assign _37 = _334;
    always @(posedge _42) begin
        if (_40)
            i_0 <= _109;
        else
            i_0 <= _37;
    end
    assign _112 = i_0 + _111;
    assign _114 = _112 == _113;
    assign _347 = _114 ? _346 : _344;
    assign _348 = _58 ? _347 : _86;
    assign _340 = _86 + _339;
    assign _342 = _88 ? _341 : _340;
    assign _338 = STATE == _63;
    assign _343 = _338 ? _342 : _86;
    assign _337 = STATE == _51;
    assign _349 = _337 ? _348 : _343;
    assign _336 = STATE == _61;
    assign _353 = _336 ? _352 : _349;
    assign _335 = STATE == _67;
    assign _356 = _335 ? _355 : _353;
    assign _38 = _356;
    always @(posedge _42) begin
        if (_40)
            _86 <= _85;
        else
            _86 <= _38;
    end
    assign _88 = _86 == _87;
    assign _372 = _88 ? _70 : STATE;
    assign _40 = clear;
    assign _42 = clock;
    assign _58 = _56 == _57;
    assign _363 = _58 ? _362 : _360;
    assign _360 = _56 + _359;
    assign _358 = STATE == _70;
    assign _361 = _358 ? _360 : _56;
    assign _357 = STATE == _51;
    assign _364 = _357 ? _363 : _361;
    assign _43 = _364;
    always @(posedge _42) begin
        if (_40)
            _56 <= _55;
        else
            _56 <= _43;
    end
    assign _76 = _56 == _75;
    assign _370 = _76 ? _67 : STATE;
    assign _369 = STATE == _70;
    assign _371 = _369 ? _370 : STATE;
    assign _368 = STATE == _63;
    assign _373 = _368 ? _372 : _371;
    assign _367 = STATE == _51;
    assign _377 = _367 ? _376 : _373;
    assign _366 = STATE == _61;
    assign _380 = _366 ? _379 : _377;
    assign _365 = STATE == _67;
    assign _382 = _365 ? _381 : _380;
    assign _44 = _382;
    always @(posedge _42) begin
        if (_40)
            STATE <= _48;
        else
            STATE <= _44;
    end
    assign _383 = STATE == _67;
    assign _398 = _383 ? _397 : _395;
    assign _45 = _398;
    always @(posedge _42) begin
        if (_40)
            _387 <= vdd;
        else
            _387 <= _45;
    end

    /* aliases */

    /* output assignments */
    assign done_ = _387;
    assign i = i_0;
    assign j = j_0;
    assign k = k_0;
    assign m = m_0;
    assign addr1 = _286;
    assign addr2 = _86;
    assign omegas0 = _280;
    assign omegas1 = _267;
    assign omegas2 = _254;
    assign omegas3 = _241;
    assign omegas4 = _228;
    assign omegas5 = _215;
    assign omegas6 = _202;
    assign start_twiddles = _189;
    assign first_stage = _148;
    assign last_stage = _128;
    assign twiddle_stage = _101;
    assign valid = _74;
    assign index = _56;
    assign read_write_enable = _3;
    assign flip = _1;

endmodule
module twdl (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    clock,
    start_twiddles,
    w
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input clock;
    input start_twiddles;
    output [63:0] w;

    /* signal declarations */
    wire [63:0] _36 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _35 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _87 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _83 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _84;
    wire [64:0] _80 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _77 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _76 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _73 = 33'b000000000000000000000000000000000;
    wire [64:0] _74;
    wire [31:0] _70 = 32'b00000000000000000000000000000000;
    wire [31:0] _69;
    wire [63:0] _71;
    wire [64:0] _72;
    wire [64:0] _75;
    reg [64:0] _78;
    wire [64:0] _67 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _66 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _63 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _61;
    wire [64:0] _62;
    wire [64:0] _64;
    wire [31:0] _57;
    wire [32:0] _56 = 33'b000000000000000000000000000000000;
    wire [64:0] _58;
    wire [127:0] _52 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _51 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _49 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _48 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _46 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _45 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _42 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _41 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _2;
    reg [63:0] _43;
    wire [63:0] _39 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    reg [63:0] _40;
    wire [127:0] _44;
    reg [127:0] _47;
    reg [127:0] _50;
    reg [127:0] _53;
    wire [63:0] _54;
    wire gnd = 1'b0;
    wire [64:0] _55;
    wire [64:0] _59;
    wire _60;
    wire [64:0] _65;
    reg [64:0] _68;
    wire [64:0] _79;
    wire _81;
    wire _82;
    wire [64:0] _85;
    wire [63:0] _86;
    reg [63:0] _89;
    wire [63:0] _4;
    wire [63:0] _6;
    wire [63:0] _8;
    wire [63:0] _10;
    wire [63:0] _12;
    wire [63:0] _14;
    wire vdd = 1'b1;
    wire [2:0] _23 = 3'b000;
    wire [2:0] _22 = 3'b000;
    wire _16;
    wire [2:0] _32 = 3'b000;
    wire [2:0] _29 = 3'b001;
    wire [2:0] _30;
    wire [2:0] _26 = 3'b110;
    wire _27;
    wire _28;
    wire [2:0] _31;
    wire [2:0] _33;
    wire [2:0] _17;
    reg [2:0] _25;
    reg [63:0] _90;
    wire _19;
    wire [63:0] _92;
    wire [63:0] _20;
    reg [63:0] _37;

    /* logic */
    assign _84 = _79 - _83;
    assign _74 = { _73, _69 };
    assign _69 = _53[95:64];
    assign _71 = { _69, _70 };
    assign _72 = { gnd, _71 };
    assign _75 = _72 - _74;
    always @(posedge _16) begin
        _78 <= _75;
    end
    assign _61 = _59[63:0];
    assign _62 = { gnd, _61 };
    assign _64 = _62 - _63;
    assign _57 = _53[127:96];
    assign _58 = { _56, _57 };
    assign _2 = omegas6;
    always @(posedge _16) begin
        _43 <= _2;
    end
    always @(posedge _16) begin
        _40 <= _37;
    end
    assign _44 = _40 * _43;
    always @(posedge _16) begin
        _47 <= _44;
    end
    always @(posedge _16) begin
        _50 <= _47;
    end
    always @(posedge _16) begin
        _53 <= _50;
    end
    assign _54 = _53[63:0];
    assign _55 = { gnd, _54 };
    assign _59 = _55 - _58;
    assign _60 = _59[64:64];
    assign _65 = _60 ? _64 : _59;
    always @(posedge _16) begin
        _68 <= _65;
    end
    assign _79 = _68 + _78;
    assign _81 = _79 < _80;
    assign _82 = ~ _81;
    assign _85 = _82 ? _84 : _79;
    assign _86 = _85[63:0];
    always @(posedge _16) begin
        _89 <= _86;
    end
    assign _4 = omegas5;
    assign _6 = omegas4;
    assign _8 = omegas3;
    assign _10 = omegas2;
    assign _12 = omegas1;
    assign _14 = omegas0;
    assign _16 = clock;
    assign _30 = _25 + _29;
    assign _27 = _25 == _26;
    assign _28 = ~ _27;
    assign _31 = _28 ? _30 : _25;
    assign _33 = _19 ? _32 : _31;
    assign _17 = _33;
    always @(posedge _16) begin
        _25 <= _17;
    end
    always @* begin
        case (_25)
        0: _90 <= _14;
        1: _90 <= _12;
        2: _90 <= _10;
        3: _90 <= _8;
        4: _90 <= _6;
        5: _90 <= _4;
        default: _90 <= _89;
        endcase
    end
    assign _19 = start_twiddles;
    assign _92 = _19 ? _91 : _90;
    assign _20 = _92;
    always @(posedge _16) begin
        _37 <= _20;
    end

    /* aliases */

    /* output assignments */
    assign w = _37;

endmodule
module dp (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_0 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0111100011111000100100011001110110001000111111001001110111000100;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0101110011101101011011100000101010001101111010000100010000101010;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1100101110010110111000101000001011011101000101101100110010111011;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0100101100101010000110001010110111100110011100100100011010110101;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0111010011110000101111011111001101001010101110111011001111101110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1110101010011101010110100001001100110110111110111100100110001011;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1000011011001101110011000011000111000011000001111110000101110001;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_1 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0000101000011000111111101100011111011101011101011111000010111001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1110100111111101110111001000100000111011101101000001000000101001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1100110100011111000010100001011101001011100011010101101111000110;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1111010100000010101011101111010100110010001100100010011001010100;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0101110011101101011011100000101010001101111010000100010000101010;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0100101100101010000110001010110111100110011100100100011010110101;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1110101010011101010110100001001100110110111110111100100110001011;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_2 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0111010000100110001111001000111100111011110010111011011011111001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1111011001111000001001110011001110101011000101110000100110010000;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0010000100100010111110011011000001011110111001100011000101100111;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1110100111111101110111001000100000111011101101000001000000101001;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1000000110000100011111010011111110001100111000110111011110101010;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0101110011101101011011100000101010001101111010000100010000101010;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0111010011110000101111011111001101001010101110111011001111101110;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_3 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0000110110101000001001111111111011110100101101110111101011101101;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0010101111111100010110000001100000101010110111101101100011110100;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1100101111011100100111001010001111010111100111010001110111111011;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0011000010111010001011101100110101011110100100111110011101101101;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1110100111111101110111001000100000111011101101000001000000101001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1111010100000010101011101111010100110010001100100010011001010100;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0100101100101010000110001010110111100110011100100100011010110101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_4 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0111110011001000110011000001001011011101111010111000111010000010;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1101100000000001010001101110001110101111011110010110111001001011;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0001011011011100101011001111000010100111110000010001101011100101;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1100101111011100100111001010001111010111100111010001110111111011;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0010000100100010111110011011000001011110111001100011000101100111;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1100110100011111000010100001011101001011100011010101101111000110;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1100101110010110111000101000001011011101000101101100110010111011;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_5 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0010101001001000011111010001011101101011111100000111111100100010;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0110110010110000111011001100000000010111101011101101100010111100;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1101100000000001010001101110001110101111011110010110111001001011;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0010101111111100010110000001100000101010110111101101100011110100;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1111011001111000001001110011001110101011000101110000100110010000;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1110100111111101110111001000100000111011101101000001000000101001;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0101110011101101011011100000101010001101111010000100010000101010;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_6 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0010100101000101111001010011010000000110010111011010001100101101;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0010101001001000011111010001011101101011111100000111111100100010;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0111110011001000110011000001001011011101111010111000111010000010;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0000110110101000001001111111111011110100101101110111101011101101;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0111010000100110001111001000111100111011110010111011011011111001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0000101000011000111111101100011111011101011101011111000010111001;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0111100011111000100100011001110110001000111111001001110111000100;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module parallel_cores (
    wr_d7,
    wr_d6,
    wr_d5,
    wr_d4,
    wr_d3,
    wr_d2,
    wr_d1,
    wr_d0,
    wr_addr,
    wr_en,
    rd_addr,
    rd_en,
    flip,
    first_4step_pass,
    first_iter,
    start,
    clear,
    clock,
    done_,
    rd_q0,
    rd_q1,
    rd_q2,
    rd_q3,
    rd_q4,
    rd_q5,
    rd_q6,
    rd_q7
);

    input [63:0] wr_d7;
    input [63:0] wr_d6;
    input [63:0] wr_d5;
    input [63:0] wr_d4;
    input [63:0] wr_d3;
    input [63:0] wr_d2;
    input [63:0] wr_d1;
    input [63:0] wr_d0;
    input [11:0] wr_addr;
    input [7:0] wr_en;
    input [11:0] rd_addr;
    input [7:0] rd_en;
    input flip;
    input first_4step_pass;
    input first_iter;
    input start;
    input clear;
    input clock;
    output done_;
    output [63:0] rd_q0;
    output [63:0] rd_q1;
    output [63:0] rd_q2;
    output [63:0] rd_q3;
    output [63:0] rd_q4;
    output [63:0] rd_q5;
    output [63:0] rd_q6;
    output [63:0] rd_q7;

    /* signal declarations */
    wire [11:0] address;
    wire write_enable;
    wire [11:0] address_0;
    wire _374;
    wire read_enable;
    wire _372;
    wire write_enable_0;
    wire _376;
    wire [131:0] _381;
    wire [63:0] _382;
    wire [11:0] _367 = 12'b000000000000;
    wire [11:0] address_1;
    wire _365;
    wire write_enable_1;
    wire [63:0] _279;
    wire [63:0] _278;
    wire [63:0] _280;
    wire [63:0] _276;
    wire [63:0] _275;
    wire [63:0] q1;
    wire [63:0] _281;
    wire [11:0] address_2;
    wire write_enable_2 = 1'b0;
    wire _266;
    wire read_enable_0;
    wire [11:0] address_3;
    wire _262;
    wire read_enable_1;
    wire _260;
    wire write_enable_3;
    wire _264;
    wire [131:0] _271;
    wire [63:0] _272;
    wire [63:0] data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_0;
    wire [11:0] _254 = 12'b000000000000;
    wire _252;
    wire _251;
    wire _250;
    wire _249;
    wire _248;
    wire _247;
    wire _246;
    wire _245;
    wire _244;
    wire _243;
    wire _242;
    wire _241;
    wire [11:0] _253;
    wire [11:0] address_4;
    wire write_enable_4 = 1'b0;
    wire _238;
    wire read_enable_2;
    wire [63:0] data_1;
    wire [63:0] data_2;
    wire _235;
    wire _234;
    wire _233;
    wire _232;
    wire _231;
    wire _230;
    wire _229;
    wire _228;
    wire _227;
    wire _226;
    wire _225;
    wire _224;
    wire [11:0] _236;
    wire [11:0] address_5;
    wire _221;
    wire read_enable_3;
    wire _219;
    wire write_enable_5;
    wire _223;
    wire [131:0] _258;
    wire [63:0] _259;
    wire _87 = 1'b0;
    wire _86 = 1'b0;
    wire _89;
    wire _3;
    reg PHASE;
    wire [63:0] _273;
    wire [11:0] address_6;
    wire _211;
    wire read_enable_4;
    wire write_enable_6;
    wire _213;
    wire [11:0] address_7;
    wire _206;
    wire read_enable_5;
    wire _204;
    wire write_enable_7;
    wire _208;
    wire [131:0] _216;
    wire [63:0] _217;
    wire [63:0] _295;
    wire [63:0] data_3;
    wire [63:0] data_4;
    wire [63:0] data_5;
    wire [63:0] data_6;
    wire [11:0] address_8;
    wire _169;
    wire read_enable_6;
    wire _166;
    wire _167;
    wire write_enable_8;
    wire _171;
    wire [11:0] address_9;
    wire _134;
    wire read_enable_7;
    wire _131;
    wire _132;
    wire write_enable_9;
    wire _136;
    wire [131:0] _202;
    wire [63:0] _203;
    wire _98 = 1'b0;
    wire _97 = 1'b0;
    wire _296;
    wire _5;
    reg PHASE_0;
    wire [63:0] q0;
    wire _94 = 1'b0;
    wire _93 = 1'b0;
    reg _96;
    wire [63:0] _274;
    wire [191:0] _294;
    wire [63:0] _297;
    wire [63:0] data_7;
    wire [63:0] data_8;
    wire [63:0] data_9;
    wire [63:0] data_10;
    wire [11:0] address_10;
    wire _361;
    wire _360;
    wire read_enable_8;
    wire _354 = 1'b0;
    wire _353 = 1'b0;
    wire _351 = 1'b0;
    wire _350 = 1'b0;
    wire _348 = 1'b0;
    wire _347 = 1'b0;
    wire _345 = 1'b0;
    wire _344 = 1'b0;
    wire _342 = 1'b0;
    wire _341 = 1'b0;
    wire _339 = 1'b0;
    wire _338 = 1'b0;
    wire _336 = 1'b0;
    wire _335 = 1'b0;
    wire _333 = 1'b0;
    wire _332 = 1'b0;
    wire _330 = 1'b0;
    wire _329 = 1'b0;
    reg _331;
    reg _334;
    reg _337;
    reg _340;
    reg _343;
    reg _346;
    reg _349;
    reg _352;
    reg _355;
    wire _356;
    wire _327 = 1'b0;
    wire _326 = 1'b0;
    wire _324 = 1'b0;
    wire _323 = 1'b0;
    wire _321 = 1'b0;
    wire _320 = 1'b0;
    wire _318 = 1'b0;
    wire _317 = 1'b0;
    wire _315 = 1'b0;
    wire _314 = 1'b0;
    wire _312 = 1'b0;
    wire _311 = 1'b0;
    wire _309 = 1'b0;
    wire _308 = 1'b0;
    wire _306 = 1'b0;
    wire _305 = 1'b0;
    wire _303 = 1'b0;
    wire _302 = 1'b0;
    reg _304;
    reg _307;
    reg _310;
    reg _313;
    reg _316;
    reg _319;
    reg _322;
    reg _325;
    reg _328;
    wire _357;
    wire _358;
    wire write_enable_10;
    wire _363;
    wire [131:0] _370;
    wire [63:0] _371;
    wire _299 = 1'b0;
    wire _298 = 1'b0;
    wire _301;
    wire _7;
    reg PHASE_1;
    wire [63:0] _383;
    wire [11:0] address_11;
    wire write_enable_11;
    wire [11:0] address_12;
    wire _570;
    wire read_enable_9;
    wire _568;
    wire write_enable_12;
    wire _572;
    wire [131:0] _577;
    wire [63:0] _578;
    wire [11:0] _563 = 12'b000000000000;
    wire [11:0] address_13;
    wire _561;
    wire write_enable_13;
    wire [63:0] _486;
    wire [63:0] _485;
    wire [63:0] _487;
    wire [63:0] _483;
    wire [63:0] _482;
    wire [63:0] q1_0;
    wire [63:0] _488;
    wire [11:0] address_14;
    wire write_enable_14 = 1'b0;
    wire _473;
    wire read_enable_10;
    wire [11:0] address_15;
    wire _469;
    wire read_enable_11;
    wire _467;
    wire write_enable_15;
    wire _471;
    wire [131:0] _478;
    wire [63:0] _479;
    wire [63:0] data_11 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_12;
    wire [11:0] _461 = 12'b000000000000;
    wire _459;
    wire _458;
    wire _457;
    wire _456;
    wire _455;
    wire _454;
    wire _453;
    wire _452;
    wire _451;
    wire _450;
    wire _449;
    wire _448;
    wire [11:0] _460;
    wire [11:0] address_16;
    wire write_enable_16 = 1'b0;
    wire _445;
    wire read_enable_12;
    wire [63:0] data_13;
    wire [63:0] data_14;
    wire _442;
    wire _441;
    wire _440;
    wire _439;
    wire _438;
    wire _437;
    wire _436;
    wire _435;
    wire _434;
    wire _433;
    wire _432;
    wire _431;
    wire [11:0] _443;
    wire [11:0] address_17;
    wire _428;
    wire read_enable_13;
    wire _426;
    wire write_enable_17;
    wire _430;
    wire [131:0] _465;
    wire [63:0] _466;
    wire _385 = 1'b0;
    wire _384 = 1'b0;
    wire _387;
    wire _11;
    reg PHASE_2;
    wire [63:0] _480;
    wire [11:0] address_18;
    wire _418;
    wire read_enable_14;
    wire write_enable_18;
    wire _420;
    wire [11:0] address_19;
    wire _413;
    wire read_enable_15;
    wire _411;
    wire write_enable_19;
    wire _415;
    wire [131:0] _423;
    wire [63:0] _424;
    wire [63:0] _491;
    wire [63:0] data_15;
    wire [63:0] data_16;
    wire [63:0] data_17;
    wire [63:0] data_18;
    wire [11:0] address_20;
    wire _404;
    wire read_enable_16;
    wire _401;
    wire _402;
    wire write_enable_20;
    wire _406;
    wire [11:0] address_21;
    wire _397;
    wire read_enable_17;
    wire _394;
    wire _395;
    wire write_enable_21;
    wire _399;
    wire [131:0] _409;
    wire [63:0] _410;
    wire _392 = 1'b0;
    wire _391 = 1'b0;
    wire _492;
    wire _13;
    reg PHASE_3;
    wire [63:0] q0_0;
    wire _389 = 1'b0;
    wire _388 = 1'b0;
    reg _390;
    wire [63:0] _481;
    wire [191:0] _490;
    wire [63:0] _493;
    wire [63:0] data_19;
    wire [63:0] data_20;
    wire [63:0] data_21;
    wire [63:0] data_22;
    wire [11:0] address_22;
    wire _557;
    wire _556;
    wire read_enable_18;
    wire _550 = 1'b0;
    wire _549 = 1'b0;
    wire _547 = 1'b0;
    wire _546 = 1'b0;
    wire _544 = 1'b0;
    wire _543 = 1'b0;
    wire _541 = 1'b0;
    wire _540 = 1'b0;
    wire _538 = 1'b0;
    wire _537 = 1'b0;
    wire _535 = 1'b0;
    wire _534 = 1'b0;
    wire _532 = 1'b0;
    wire _531 = 1'b0;
    wire _529 = 1'b0;
    wire _528 = 1'b0;
    wire _526 = 1'b0;
    wire _525 = 1'b0;
    reg _527;
    reg _530;
    reg _533;
    reg _536;
    reg _539;
    reg _542;
    reg _545;
    reg _548;
    reg _551;
    wire _552;
    wire _523 = 1'b0;
    wire _522 = 1'b0;
    wire _520 = 1'b0;
    wire _519 = 1'b0;
    wire _517 = 1'b0;
    wire _516 = 1'b0;
    wire _514 = 1'b0;
    wire _513 = 1'b0;
    wire _511 = 1'b0;
    wire _510 = 1'b0;
    wire _508 = 1'b0;
    wire _507 = 1'b0;
    wire _505 = 1'b0;
    wire _504 = 1'b0;
    wire _502 = 1'b0;
    wire _501 = 1'b0;
    wire _499 = 1'b0;
    wire _498 = 1'b0;
    reg _500;
    reg _503;
    reg _506;
    reg _509;
    reg _512;
    reg _515;
    reg _518;
    reg _521;
    reg _524;
    wire _553;
    wire _554;
    wire write_enable_22;
    wire _559;
    wire [131:0] _566;
    wire [63:0] _567;
    wire _495 = 1'b0;
    wire _494 = 1'b0;
    wire _497;
    wire _15;
    reg PHASE_4;
    wire [63:0] _579;
    wire [11:0] address_23;
    wire write_enable_23;
    wire [11:0] address_24;
    wire _766;
    wire read_enable_19;
    wire _764;
    wire write_enable_24;
    wire _768;
    wire [131:0] _773;
    wire [63:0] _774;
    wire [11:0] _759 = 12'b000000000000;
    wire [11:0] address_25;
    wire _757;
    wire write_enable_25;
    wire [63:0] _682;
    wire [63:0] _681;
    wire [63:0] _683;
    wire [63:0] _679;
    wire [63:0] _678;
    wire [63:0] q1_1;
    wire [63:0] _684;
    wire [11:0] address_26;
    wire write_enable_26 = 1'b0;
    wire _669;
    wire read_enable_20;
    wire [11:0] address_27;
    wire _665;
    wire read_enable_21;
    wire _663;
    wire write_enable_27;
    wire _667;
    wire [131:0] _674;
    wire [63:0] _675;
    wire [63:0] data_23 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_24;
    wire [11:0] _657 = 12'b000000000000;
    wire _655;
    wire _654;
    wire _653;
    wire _652;
    wire _651;
    wire _650;
    wire _649;
    wire _648;
    wire _647;
    wire _646;
    wire _645;
    wire _644;
    wire [11:0] _656;
    wire [11:0] address_28;
    wire write_enable_28 = 1'b0;
    wire _641;
    wire read_enable_22;
    wire [63:0] data_25;
    wire [63:0] data_26;
    wire _638;
    wire _637;
    wire _636;
    wire _635;
    wire _634;
    wire _633;
    wire _632;
    wire _631;
    wire _630;
    wire _629;
    wire _628;
    wire _627;
    wire [11:0] _639;
    wire [11:0] address_29;
    wire _624;
    wire read_enable_23;
    wire _622;
    wire write_enable_29;
    wire _626;
    wire [131:0] _661;
    wire [63:0] _662;
    wire _581 = 1'b0;
    wire _580 = 1'b0;
    wire _583;
    wire _19;
    reg PHASE_5;
    wire [63:0] _676;
    wire [11:0] address_30;
    wire _614;
    wire read_enable_24;
    wire write_enable_30;
    wire _616;
    wire [11:0] address_31;
    wire _609;
    wire read_enable_25;
    wire _607;
    wire write_enable_31;
    wire _611;
    wire [131:0] _619;
    wire [63:0] _620;
    wire [63:0] _687;
    wire [63:0] data_27;
    wire [63:0] data_28;
    wire [63:0] data_29;
    wire [63:0] data_30;
    wire [11:0] address_32;
    wire _600;
    wire read_enable_26;
    wire _597;
    wire _598;
    wire write_enable_32;
    wire _602;
    wire [11:0] address_33;
    wire _593;
    wire read_enable_27;
    wire _590;
    wire _591;
    wire write_enable_33;
    wire _595;
    wire [131:0] _605;
    wire [63:0] _606;
    wire _588 = 1'b0;
    wire _587 = 1'b0;
    wire _688;
    wire _21;
    reg PHASE_6;
    wire [63:0] q0_1;
    wire _585 = 1'b0;
    wire _584 = 1'b0;
    reg _586;
    wire [63:0] _677;
    wire [191:0] _686;
    wire [63:0] _689;
    wire [63:0] data_31;
    wire [63:0] data_32;
    wire [63:0] data_33;
    wire [63:0] data_34;
    wire [11:0] address_34;
    wire _753;
    wire _752;
    wire read_enable_28;
    wire _746 = 1'b0;
    wire _745 = 1'b0;
    wire _743 = 1'b0;
    wire _742 = 1'b0;
    wire _740 = 1'b0;
    wire _739 = 1'b0;
    wire _737 = 1'b0;
    wire _736 = 1'b0;
    wire _734 = 1'b0;
    wire _733 = 1'b0;
    wire _731 = 1'b0;
    wire _730 = 1'b0;
    wire _728 = 1'b0;
    wire _727 = 1'b0;
    wire _725 = 1'b0;
    wire _724 = 1'b0;
    wire _722 = 1'b0;
    wire _721 = 1'b0;
    reg _723;
    reg _726;
    reg _729;
    reg _732;
    reg _735;
    reg _738;
    reg _741;
    reg _744;
    reg _747;
    wire _748;
    wire _719 = 1'b0;
    wire _718 = 1'b0;
    wire _716 = 1'b0;
    wire _715 = 1'b0;
    wire _713 = 1'b0;
    wire _712 = 1'b0;
    wire _710 = 1'b0;
    wire _709 = 1'b0;
    wire _707 = 1'b0;
    wire _706 = 1'b0;
    wire _704 = 1'b0;
    wire _703 = 1'b0;
    wire _701 = 1'b0;
    wire _700 = 1'b0;
    wire _698 = 1'b0;
    wire _697 = 1'b0;
    wire _695 = 1'b0;
    wire _694 = 1'b0;
    reg _696;
    reg _699;
    reg _702;
    reg _705;
    reg _708;
    reg _711;
    reg _714;
    reg _717;
    reg _720;
    wire _749;
    wire _750;
    wire write_enable_34;
    wire _755;
    wire [131:0] _762;
    wire [63:0] _763;
    wire _691 = 1'b0;
    wire _690 = 1'b0;
    wire _693;
    wire _23;
    reg PHASE_7;
    wire [63:0] _775;
    wire [11:0] address_35;
    wire write_enable_35;
    wire [11:0] address_36;
    wire _962;
    wire read_enable_29;
    wire _960;
    wire write_enable_36;
    wire _964;
    wire [131:0] _969;
    wire [63:0] _970;
    wire [11:0] _955 = 12'b000000000000;
    wire [11:0] address_37;
    wire _953;
    wire write_enable_37;
    wire [63:0] _878;
    wire [63:0] _877;
    wire [63:0] _879;
    wire [63:0] _875;
    wire [63:0] _874;
    wire [63:0] q1_2;
    wire [63:0] _880;
    wire [11:0] address_38;
    wire write_enable_38 = 1'b0;
    wire _865;
    wire read_enable_30;
    wire [11:0] address_39;
    wire _861;
    wire read_enable_31;
    wire _859;
    wire write_enable_39;
    wire _863;
    wire [131:0] _870;
    wire [63:0] _871;
    wire [63:0] data_35 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_36;
    wire [11:0] _853 = 12'b000000000000;
    wire _851;
    wire _850;
    wire _849;
    wire _848;
    wire _847;
    wire _846;
    wire _845;
    wire _844;
    wire _843;
    wire _842;
    wire _841;
    wire _840;
    wire [11:0] _852;
    wire [11:0] address_40;
    wire write_enable_40 = 1'b0;
    wire _837;
    wire read_enable_32;
    wire [63:0] data_37;
    wire [63:0] data_38;
    wire _834;
    wire _833;
    wire _832;
    wire _831;
    wire _830;
    wire _829;
    wire _828;
    wire _827;
    wire _826;
    wire _825;
    wire _824;
    wire _823;
    wire [11:0] _835;
    wire [11:0] address_41;
    wire _820;
    wire read_enable_33;
    wire _818;
    wire write_enable_41;
    wire _822;
    wire [131:0] _857;
    wire [63:0] _858;
    wire _777 = 1'b0;
    wire _776 = 1'b0;
    wire _779;
    wire _27;
    reg PHASE_8;
    wire [63:0] _872;
    wire [11:0] address_42;
    wire _810;
    wire read_enable_34;
    wire write_enable_42;
    wire _812;
    wire [11:0] address_43;
    wire _805;
    wire read_enable_35;
    wire _803;
    wire write_enable_43;
    wire _807;
    wire [131:0] _815;
    wire [63:0] _816;
    wire [63:0] _883;
    wire [63:0] data_39;
    wire [63:0] data_40;
    wire [63:0] data_41;
    wire [63:0] data_42;
    wire [11:0] address_44;
    wire _796;
    wire read_enable_36;
    wire _793;
    wire _794;
    wire write_enable_44;
    wire _798;
    wire [11:0] address_45;
    wire _789;
    wire read_enable_37;
    wire _786;
    wire _787;
    wire write_enable_45;
    wire _791;
    wire [131:0] _801;
    wire [63:0] _802;
    wire _784 = 1'b0;
    wire _783 = 1'b0;
    wire _884;
    wire _29;
    reg PHASE_9;
    wire [63:0] q0_2;
    wire _781 = 1'b0;
    wire _780 = 1'b0;
    reg _782;
    wire [63:0] _873;
    wire [191:0] _882;
    wire [63:0] _885;
    wire [63:0] data_43;
    wire [63:0] data_44;
    wire [63:0] data_45;
    wire [63:0] data_46;
    wire [11:0] address_46;
    wire _949;
    wire _948;
    wire read_enable_38;
    wire _942 = 1'b0;
    wire _941 = 1'b0;
    wire _939 = 1'b0;
    wire _938 = 1'b0;
    wire _936 = 1'b0;
    wire _935 = 1'b0;
    wire _933 = 1'b0;
    wire _932 = 1'b0;
    wire _930 = 1'b0;
    wire _929 = 1'b0;
    wire _927 = 1'b0;
    wire _926 = 1'b0;
    wire _924 = 1'b0;
    wire _923 = 1'b0;
    wire _921 = 1'b0;
    wire _920 = 1'b0;
    wire _918 = 1'b0;
    wire _917 = 1'b0;
    reg _919;
    reg _922;
    reg _925;
    reg _928;
    reg _931;
    reg _934;
    reg _937;
    reg _940;
    reg _943;
    wire _944;
    wire _915 = 1'b0;
    wire _914 = 1'b0;
    wire _912 = 1'b0;
    wire _911 = 1'b0;
    wire _909 = 1'b0;
    wire _908 = 1'b0;
    wire _906 = 1'b0;
    wire _905 = 1'b0;
    wire _903 = 1'b0;
    wire _902 = 1'b0;
    wire _900 = 1'b0;
    wire _899 = 1'b0;
    wire _897 = 1'b0;
    wire _896 = 1'b0;
    wire _894 = 1'b0;
    wire _893 = 1'b0;
    wire _891 = 1'b0;
    wire _890 = 1'b0;
    reg _892;
    reg _895;
    reg _898;
    reg _901;
    reg _904;
    reg _907;
    reg _910;
    reg _913;
    reg _916;
    wire _945;
    wire _946;
    wire write_enable_46;
    wire _951;
    wire [131:0] _958;
    wire [63:0] _959;
    wire _887 = 1'b0;
    wire _886 = 1'b0;
    wire _889;
    wire _31;
    reg PHASE_10;
    wire [63:0] _971;
    wire [11:0] address_47;
    wire write_enable_47;
    wire [11:0] address_48;
    wire _1158;
    wire read_enable_39;
    wire _1156;
    wire write_enable_48;
    wire _1160;
    wire [131:0] _1165;
    wire [63:0] _1166;
    wire [11:0] _1151 = 12'b000000000000;
    wire [11:0] address_49;
    wire _1149;
    wire write_enable_49;
    wire [63:0] _1074;
    wire [63:0] _1073;
    wire [63:0] _1075;
    wire [63:0] _1071;
    wire [63:0] _1070;
    wire [63:0] q1_3;
    wire [63:0] _1076;
    wire [11:0] address_50;
    wire write_enable_50 = 1'b0;
    wire _1061;
    wire read_enable_40;
    wire [11:0] address_51;
    wire _1057;
    wire read_enable_41;
    wire _1055;
    wire write_enable_51;
    wire _1059;
    wire [131:0] _1066;
    wire [63:0] _1067;
    wire [63:0] data_47 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_48;
    wire [11:0] _1049 = 12'b000000000000;
    wire _1047;
    wire _1046;
    wire _1045;
    wire _1044;
    wire _1043;
    wire _1042;
    wire _1041;
    wire _1040;
    wire _1039;
    wire _1038;
    wire _1037;
    wire _1036;
    wire [11:0] _1048;
    wire [11:0] address_52;
    wire write_enable_52 = 1'b0;
    wire _1033;
    wire read_enable_42;
    wire [63:0] data_49;
    wire [63:0] data_50;
    wire _1030;
    wire _1029;
    wire _1028;
    wire _1027;
    wire _1026;
    wire _1025;
    wire _1024;
    wire _1023;
    wire _1022;
    wire _1021;
    wire _1020;
    wire _1019;
    wire [11:0] _1031;
    wire [11:0] address_53;
    wire _1016;
    wire read_enable_43;
    wire _1014;
    wire write_enable_53;
    wire _1018;
    wire [131:0] _1053;
    wire [63:0] _1054;
    wire _973 = 1'b0;
    wire _972 = 1'b0;
    wire _975;
    wire _35;
    reg PHASE_11;
    wire [63:0] _1068;
    wire [11:0] address_54;
    wire _1006;
    wire read_enable_44;
    wire write_enable_54;
    wire _1008;
    wire [11:0] address_55;
    wire _1001;
    wire read_enable_45;
    wire _999;
    wire write_enable_55;
    wire _1003;
    wire [131:0] _1011;
    wire [63:0] _1012;
    wire [63:0] _1079;
    wire [63:0] data_51;
    wire [63:0] data_52;
    wire [63:0] data_53;
    wire [63:0] data_54;
    wire [11:0] address_56;
    wire _992;
    wire read_enable_46;
    wire _989;
    wire _990;
    wire write_enable_56;
    wire _994;
    wire [11:0] address_57;
    wire _985;
    wire read_enable_47;
    wire _982;
    wire _983;
    wire write_enable_57;
    wire _987;
    wire [131:0] _997;
    wire [63:0] _998;
    wire _980 = 1'b0;
    wire _979 = 1'b0;
    wire _1080;
    wire _37;
    reg PHASE_12;
    wire [63:0] q0_3;
    wire _977 = 1'b0;
    wire _976 = 1'b0;
    reg _978;
    wire [63:0] _1069;
    wire [191:0] _1078;
    wire [63:0] _1081;
    wire [63:0] data_55;
    wire [63:0] data_56;
    wire [63:0] data_57;
    wire [63:0] data_58;
    wire [11:0] address_58;
    wire _1145;
    wire _1144;
    wire read_enable_48;
    wire _1138 = 1'b0;
    wire _1137 = 1'b0;
    wire _1135 = 1'b0;
    wire _1134 = 1'b0;
    wire _1132 = 1'b0;
    wire _1131 = 1'b0;
    wire _1129 = 1'b0;
    wire _1128 = 1'b0;
    wire _1126 = 1'b0;
    wire _1125 = 1'b0;
    wire _1123 = 1'b0;
    wire _1122 = 1'b0;
    wire _1120 = 1'b0;
    wire _1119 = 1'b0;
    wire _1117 = 1'b0;
    wire _1116 = 1'b0;
    wire _1114 = 1'b0;
    wire _1113 = 1'b0;
    reg _1115;
    reg _1118;
    reg _1121;
    reg _1124;
    reg _1127;
    reg _1130;
    reg _1133;
    reg _1136;
    reg _1139;
    wire _1140;
    wire _1111 = 1'b0;
    wire _1110 = 1'b0;
    wire _1108 = 1'b0;
    wire _1107 = 1'b0;
    wire _1105 = 1'b0;
    wire _1104 = 1'b0;
    wire _1102 = 1'b0;
    wire _1101 = 1'b0;
    wire _1099 = 1'b0;
    wire _1098 = 1'b0;
    wire _1096 = 1'b0;
    wire _1095 = 1'b0;
    wire _1093 = 1'b0;
    wire _1092 = 1'b0;
    wire _1090 = 1'b0;
    wire _1089 = 1'b0;
    wire _1087 = 1'b0;
    wire _1086 = 1'b0;
    reg _1088;
    reg _1091;
    reg _1094;
    reg _1097;
    reg _1100;
    reg _1103;
    reg _1106;
    reg _1109;
    reg _1112;
    wire _1141;
    wire _1142;
    wire write_enable_58;
    wire _1147;
    wire [131:0] _1154;
    wire [63:0] _1155;
    wire _1083 = 1'b0;
    wire _1082 = 1'b0;
    wire _1085;
    wire _39;
    reg PHASE_13;
    wire [63:0] _1167;
    wire [11:0] address_59;
    wire write_enable_59;
    wire [11:0] address_60;
    wire _1354;
    wire read_enable_49;
    wire _1352;
    wire write_enable_60;
    wire _1356;
    wire [131:0] _1361;
    wire [63:0] _1362;
    wire [11:0] _1347 = 12'b000000000000;
    wire [11:0] address_61;
    wire _1345;
    wire write_enable_61;
    wire [63:0] _1270;
    wire [63:0] _1269;
    wire [63:0] _1271;
    wire [63:0] _1267;
    wire [63:0] _1266;
    wire [63:0] q1_4;
    wire [63:0] _1272;
    wire [11:0] address_62;
    wire write_enable_62 = 1'b0;
    wire _1257;
    wire read_enable_50;
    wire [11:0] address_63;
    wire _1253;
    wire read_enable_51;
    wire _1251;
    wire write_enable_63;
    wire _1255;
    wire [131:0] _1262;
    wire [63:0] _1263;
    wire [63:0] data_59 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_60;
    wire [11:0] _1245 = 12'b000000000000;
    wire _1243;
    wire _1242;
    wire _1241;
    wire _1240;
    wire _1239;
    wire _1238;
    wire _1237;
    wire _1236;
    wire _1235;
    wire _1234;
    wire _1233;
    wire _1232;
    wire [11:0] _1244;
    wire [11:0] address_64;
    wire write_enable_64 = 1'b0;
    wire _1229;
    wire read_enable_52;
    wire [63:0] data_61;
    wire [63:0] data_62;
    wire _1226;
    wire _1225;
    wire _1224;
    wire _1223;
    wire _1222;
    wire _1221;
    wire _1220;
    wire _1219;
    wire _1218;
    wire _1217;
    wire _1216;
    wire _1215;
    wire [11:0] _1227;
    wire [11:0] address_65;
    wire _1212;
    wire read_enable_53;
    wire _1210;
    wire write_enable_65;
    wire _1214;
    wire [131:0] _1249;
    wire [63:0] _1250;
    wire _1169 = 1'b0;
    wire _1168 = 1'b0;
    wire _1171;
    wire _43;
    reg PHASE_14;
    wire [63:0] _1264;
    wire [11:0] address_66;
    wire _1202;
    wire read_enable_54;
    wire write_enable_66;
    wire _1204;
    wire [11:0] address_67;
    wire _1197;
    wire read_enable_55;
    wire _1195;
    wire write_enable_67;
    wire _1199;
    wire [131:0] _1207;
    wire [63:0] _1208;
    wire [63:0] _1275;
    wire [63:0] data_63;
    wire [63:0] data_64;
    wire [63:0] data_65;
    wire [63:0] data_66;
    wire [11:0] address_68;
    wire _1188;
    wire read_enable_56;
    wire _1185;
    wire _1186;
    wire write_enable_68;
    wire _1190;
    wire [11:0] address_69;
    wire _1181;
    wire read_enable_57;
    wire _1178;
    wire _1179;
    wire write_enable_69;
    wire _1183;
    wire [131:0] _1193;
    wire [63:0] _1194;
    wire _1176 = 1'b0;
    wire _1175 = 1'b0;
    wire _1276;
    wire _45;
    reg PHASE_15;
    wire [63:0] q0_4;
    wire _1173 = 1'b0;
    wire _1172 = 1'b0;
    reg _1174;
    wire [63:0] _1265;
    wire [191:0] _1274;
    wire [63:0] _1277;
    wire [63:0] data_67;
    wire [63:0] data_68;
    wire [63:0] data_69;
    wire [63:0] data_70;
    wire [11:0] address_70;
    wire _1341;
    wire _1340;
    wire read_enable_58;
    wire _1334 = 1'b0;
    wire _1333 = 1'b0;
    wire _1331 = 1'b0;
    wire _1330 = 1'b0;
    wire _1328 = 1'b0;
    wire _1327 = 1'b0;
    wire _1325 = 1'b0;
    wire _1324 = 1'b0;
    wire _1322 = 1'b0;
    wire _1321 = 1'b0;
    wire _1319 = 1'b0;
    wire _1318 = 1'b0;
    wire _1316 = 1'b0;
    wire _1315 = 1'b0;
    wire _1313 = 1'b0;
    wire _1312 = 1'b0;
    wire _1310 = 1'b0;
    wire _1309 = 1'b0;
    reg _1311;
    reg _1314;
    reg _1317;
    reg _1320;
    reg _1323;
    reg _1326;
    reg _1329;
    reg _1332;
    reg _1335;
    wire _1336;
    wire _1307 = 1'b0;
    wire _1306 = 1'b0;
    wire _1304 = 1'b0;
    wire _1303 = 1'b0;
    wire _1301 = 1'b0;
    wire _1300 = 1'b0;
    wire _1298 = 1'b0;
    wire _1297 = 1'b0;
    wire _1295 = 1'b0;
    wire _1294 = 1'b0;
    wire _1292 = 1'b0;
    wire _1291 = 1'b0;
    wire _1289 = 1'b0;
    wire _1288 = 1'b0;
    wire _1286 = 1'b0;
    wire _1285 = 1'b0;
    wire _1283 = 1'b0;
    wire _1282 = 1'b0;
    reg _1284;
    reg _1287;
    reg _1290;
    reg _1293;
    reg _1296;
    reg _1299;
    reg _1302;
    reg _1305;
    reg _1308;
    wire _1337;
    wire _1338;
    wire write_enable_70;
    wire _1343;
    wire [131:0] _1350;
    wire [63:0] _1351;
    wire _1279 = 1'b0;
    wire _1278 = 1'b0;
    wire _1281;
    wire _47;
    reg PHASE_16;
    wire [63:0] _1363;
    wire [11:0] address_71;
    wire write_enable_71;
    wire [11:0] address_72;
    wire _1550;
    wire read_enable_59;
    wire _1548;
    wire write_enable_72;
    wire _1552;
    wire [131:0] _1557;
    wire [63:0] _1558;
    wire [11:0] _1543 = 12'b000000000000;
    wire [11:0] address_73;
    wire _1541;
    wire write_enable_73;
    wire [63:0] _1466;
    wire [63:0] _1465;
    wire [63:0] _1467;
    wire [63:0] _1463;
    wire [63:0] _1462;
    wire [63:0] q1_5;
    wire [63:0] _1468;
    wire [11:0] address_74;
    wire write_enable_74 = 1'b0;
    wire _1453;
    wire read_enable_60;
    wire [11:0] address_75;
    wire _1449;
    wire read_enable_61;
    wire _1447;
    wire write_enable_75;
    wire _1451;
    wire [131:0] _1458;
    wire [63:0] _1459;
    wire [63:0] data_71 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_72;
    wire [11:0] _1441 = 12'b000000000000;
    wire _1439;
    wire _1438;
    wire _1437;
    wire _1436;
    wire _1435;
    wire _1434;
    wire _1433;
    wire _1432;
    wire _1431;
    wire _1430;
    wire _1429;
    wire _1428;
    wire [11:0] _1440;
    wire [11:0] address_76;
    wire write_enable_76 = 1'b0;
    wire _1425;
    wire read_enable_62;
    wire [63:0] data_73;
    wire [63:0] data_74;
    wire _1422;
    wire _1421;
    wire _1420;
    wire _1419;
    wire _1418;
    wire _1417;
    wire _1416;
    wire _1415;
    wire _1414;
    wire _1413;
    wire _1412;
    wire _1411;
    wire [11:0] _1423;
    wire [11:0] address_77;
    wire _1408;
    wire read_enable_63;
    wire _1406;
    wire write_enable_77;
    wire _1410;
    wire [131:0] _1445;
    wire [63:0] _1446;
    wire _1365 = 1'b0;
    wire _1364 = 1'b0;
    wire _1367;
    wire _51;
    reg PHASE_17;
    wire [63:0] _1460;
    wire [11:0] address_78;
    wire _1398;
    wire read_enable_64;
    wire write_enable_78;
    wire _1400;
    wire [11:0] address_79;
    wire _1393;
    wire read_enable_65;
    wire _1391;
    wire write_enable_79;
    wire _1395;
    wire [131:0] _1403;
    wire [63:0] _1404;
    wire [63:0] _1471;
    wire [63:0] data_75;
    wire [63:0] data_76;
    wire [63:0] data_77;
    wire [63:0] data_78;
    wire [11:0] address_80;
    wire _1384;
    wire read_enable_66;
    wire _1381;
    wire _1382;
    wire write_enable_80;
    wire _1386;
    wire [11:0] address_81;
    wire _1377;
    wire read_enable_67;
    wire _1374;
    wire _1375;
    wire write_enable_81;
    wire _1379;
    wire [131:0] _1389;
    wire [63:0] _1390;
    wire _1372 = 1'b0;
    wire _1371 = 1'b0;
    wire _1472;
    wire _53;
    reg PHASE_18;
    wire [63:0] q0_5;
    wire _1369 = 1'b0;
    wire _1368 = 1'b0;
    reg _1370;
    wire [63:0] _1461;
    wire [191:0] _1470;
    wire [63:0] _1473;
    wire [63:0] data_79;
    wire [63:0] data_80;
    wire [63:0] data_81;
    wire [63:0] data_82;
    wire [11:0] address_82;
    wire _1537;
    wire _1536;
    wire read_enable_68;
    wire _1530 = 1'b0;
    wire _1529 = 1'b0;
    wire _1527 = 1'b0;
    wire _1526 = 1'b0;
    wire _1524 = 1'b0;
    wire _1523 = 1'b0;
    wire _1521 = 1'b0;
    wire _1520 = 1'b0;
    wire _1518 = 1'b0;
    wire _1517 = 1'b0;
    wire _1515 = 1'b0;
    wire _1514 = 1'b0;
    wire _1512 = 1'b0;
    wire _1511 = 1'b0;
    wire _1509 = 1'b0;
    wire _1508 = 1'b0;
    wire _1506 = 1'b0;
    wire _1505 = 1'b0;
    reg _1507;
    reg _1510;
    reg _1513;
    reg _1516;
    reg _1519;
    reg _1522;
    reg _1525;
    reg _1528;
    reg _1531;
    wire _1532;
    wire _1503 = 1'b0;
    wire _1502 = 1'b0;
    wire _1500 = 1'b0;
    wire _1499 = 1'b0;
    wire _1497 = 1'b0;
    wire _1496 = 1'b0;
    wire _1494 = 1'b0;
    wire _1493 = 1'b0;
    wire _1491 = 1'b0;
    wire _1490 = 1'b0;
    wire _1488 = 1'b0;
    wire _1487 = 1'b0;
    wire _1485 = 1'b0;
    wire _1484 = 1'b0;
    wire _1482 = 1'b0;
    wire _1481 = 1'b0;
    wire _1479 = 1'b0;
    wire _1478 = 1'b0;
    reg _1480;
    reg _1483;
    reg _1486;
    reg _1489;
    reg _1492;
    reg _1495;
    reg _1498;
    reg _1501;
    reg _1504;
    wire _1533;
    wire _1534;
    wire write_enable_82;
    wire _1539;
    wire [131:0] _1546;
    wire [63:0] _1547;
    wire _1475 = 1'b0;
    wire _1474 = 1'b0;
    wire _1477;
    wire _55;
    reg PHASE_19;
    wire [63:0] _1559;
    wire [11:0] address_83;
    wire write_enable_83;
    wire [11:0] address_84;
    wire _1746;
    wire read_enable_69;
    wire _1744;
    wire write_enable_84;
    wire _1748;
    wire [131:0] _1753;
    wire [63:0] _1754;
    wire [11:0] _1739 = 12'b000000000000;
    wire [11:0] address_85;
    wire _1737;
    wire write_enable_85;
    wire [3:0] _292;
    wire _291;
    wire _289;
    wire [63:0] _288;
    wire [63:0] _287;
    wire [63:0] _286;
    wire [63:0] _285;
    wire [63:0] _284;
    wire [63:0] _283;
    wire [63:0] _282;
    wire [63:0] _1662;
    wire [63:0] _1661;
    wire [63:0] _1663;
    wire [63:0] _1659;
    wire [63:0] _1658;
    wire [63:0] q1_6;
    wire [63:0] _1664;
    wire [11:0] address_86;
    wire write_enable_86 = 1'b0;
    wire _1649;
    wire read_enable_70;
    wire [11:0] address_87;
    wire _1645;
    wire read_enable_71;
    wire _1643;
    wire write_enable_87;
    wire _1647;
    wire [131:0] _1654;
    wire [63:0] _1655;
    wire [63:0] data_83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_84;
    wire [11:0] _1637 = 12'b000000000000;
    wire _1635;
    wire _1634;
    wire _1633;
    wire _1632;
    wire _1631;
    wire _1630;
    wire _1629;
    wire _1628;
    wire _1627;
    wire _1626;
    wire _1625;
    wire _1624;
    wire [11:0] _1636;
    wire [11:0] address_88;
    wire write_enable_88 = 1'b0;
    wire _1621;
    wire read_enable_72;
    wire [63:0] data_85;
    wire [63:0] data_86;
    wire [11:0] _60;
    wire _1618;
    wire _1617;
    wire _1616;
    wire _1615;
    wire _1614;
    wire _1613;
    wire _1612;
    wire _1611;
    wire _1610;
    wire _1609;
    wire _1608;
    wire _1607;
    wire [11:0] _1619;
    wire [11:0] address_89;
    wire _1604;
    wire read_enable_73;
    wire [7:0] _62;
    wire _1602;
    wire write_enable_89;
    wire _1606;
    wire [131:0] _1641;
    wire [63:0] _1642;
    wire _1561 = 1'b0;
    wire _1560 = 1'b0;
    wire _1563;
    wire _63;
    reg PHASE_20;
    wire [63:0] _1656;
    wire [11:0] address_90;
    wire _1594;
    wire read_enable_74;
    wire write_enable_90;
    wire _1596;
    wire [11:0] address_91;
    wire _1589;
    wire read_enable_75;
    wire _1587;
    wire write_enable_91;
    wire _1591;
    wire [131:0] _1599;
    wire [63:0] _1600;
    wire [63:0] _1667;
    wire [63:0] data_87;
    wire [63:0] data_88;
    wire [63:0] data_89;
    wire [63:0] data_90;
    wire [11:0] _198 = 12'b000000000000;
    wire [11:0] _197 = 12'b000000000000;
    wire [11:0] _195 = 12'b000000000000;
    wire [11:0] _194 = 12'b000000000000;
    wire [11:0] _192 = 12'b000000000000;
    wire [11:0] _191 = 12'b000000000000;
    wire [11:0] _189 = 12'b000000000000;
    wire [11:0] _188 = 12'b000000000000;
    wire [11:0] _186 = 12'b000000000000;
    wire [11:0] _185 = 12'b000000000000;
    wire [11:0] _183 = 12'b000000000000;
    wire [11:0] _182 = 12'b000000000000;
    wire [11:0] _180 = 12'b000000000000;
    wire [11:0] _179 = 12'b000000000000;
    wire [11:0] _177 = 12'b000000000000;
    wire [11:0] _176 = 12'b000000000000;
    wire [11:0] _174 = 12'b000000000000;
    wire [11:0] _173 = 12'b000000000000;
    reg [11:0] _175;
    reg [11:0] _178;
    reg [11:0] _181;
    reg [11:0] _184;
    reg [11:0] _187;
    reg [11:0] _190;
    reg [11:0] _193;
    reg [11:0] _196;
    reg [11:0] _199;
    wire [11:0] _172;
    wire [11:0] address_92;
    wire _1580;
    wire read_enable_76;
    wire _1577;
    wire _1578;
    wire write_enable_92;
    wire _1582;
    wire [11:0] address_93;
    wire _1573;
    wire read_enable_77;
    wire _1570;
    wire _1571;
    wire write_enable_93;
    wire _1575;
    wire [131:0] _1585;
    wire [63:0] _1586;
    wire _99;
    wire _1568 = 1'b0;
    wire _1567 = 1'b0;
    wire _1668;
    wire _65;
    reg PHASE_21;
    wire [63:0] q0_6;
    wire _1565 = 1'b0;
    wire _1564 = 1'b0;
    wire _92;
    reg _1566;
    wire [63:0] _1657;
    wire [191:0] _1666;
    wire [63:0] _1669;
    wire [63:0] data_91;
    wire [63:0] data_92;
    wire [63:0] data_93;
    wire [63:0] data_94;
    wire [11:0] _163 = 12'b000000000000;
    wire [11:0] _162 = 12'b000000000000;
    wire [11:0] _160 = 12'b000000000000;
    wire [11:0] _159 = 12'b000000000000;
    wire [11:0] _157 = 12'b000000000000;
    wire [11:0] _156 = 12'b000000000000;
    wire [11:0] _154 = 12'b000000000000;
    wire [11:0] _153 = 12'b000000000000;
    wire [11:0] _151 = 12'b000000000000;
    wire [11:0] _150 = 12'b000000000000;
    wire [11:0] _148 = 12'b000000000000;
    wire [11:0] _147 = 12'b000000000000;
    wire [11:0] _145 = 12'b000000000000;
    wire [11:0] _144 = 12'b000000000000;
    wire [11:0] _142 = 12'b000000000000;
    wire [11:0] _141 = 12'b000000000000;
    wire [11:0] _139 = 12'b000000000000;
    wire [11:0] _138 = 12'b000000000000;
    wire [11:0] _137;
    reg [11:0] _140;
    reg [11:0] _143;
    reg [11:0] _146;
    reg [11:0] _149;
    reg [11:0] _152;
    reg [11:0] _155;
    reg [11:0] _158;
    reg [11:0] _161;
    reg [11:0] _164;
    wire [11:0] _68;
    wire [11:0] address_94;
    wire _1733;
    wire [7:0] _70;
    wire _1732;
    wire read_enable_78;
    wire _1726 = 1'b0;
    wire _1725 = 1'b0;
    wire _1723 = 1'b0;
    wire _1722 = 1'b0;
    wire _1720 = 1'b0;
    wire _1719 = 1'b0;
    wire _1717 = 1'b0;
    wire _1716 = 1'b0;
    wire _1714 = 1'b0;
    wire _1713 = 1'b0;
    wire _1711 = 1'b0;
    wire _1710 = 1'b0;
    wire _1708 = 1'b0;
    wire _1707 = 1'b0;
    wire _1705 = 1'b0;
    wire _1704 = 1'b0;
    wire _1702 = 1'b0;
    wire _1701 = 1'b0;
    wire _290;
    reg _1703;
    reg _1706;
    reg _1709;
    reg _1712;
    reg _1715;
    reg _1718;
    reg _1721;
    reg _1724;
    reg _1727;
    wire _1728;
    wire _1699 = 1'b0;
    wire _1698 = 1'b0;
    wire _1696 = 1'b0;
    wire _1695 = 1'b0;
    wire _1693 = 1'b0;
    wire _1692 = 1'b0;
    wire _1690 = 1'b0;
    wire _1689 = 1'b0;
    wire _1687 = 1'b0;
    wire _1686 = 1'b0;
    wire _1684 = 1'b0;
    wire _1683 = 1'b0;
    wire _1681 = 1'b0;
    wire _1680 = 1'b0;
    wire _1678 = 1'b0;
    wire _1677 = 1'b0;
    wire _1675 = 1'b0;
    wire _1674 = 1'b0;
    wire _130;
    reg _1676;
    reg _1679;
    reg _1682;
    reg _1685;
    reg _1688;
    reg _1691;
    reg _1694;
    reg _1697;
    reg _1700;
    wire _1729;
    wire _128 = 1'b0;
    wire _127 = 1'b0;
    wire _125 = 1'b0;
    wire _124 = 1'b0;
    wire _122 = 1'b0;
    wire _121 = 1'b0;
    wire _119 = 1'b0;
    wire _118 = 1'b0;
    wire _116 = 1'b0;
    wire _115 = 1'b0;
    wire _113 = 1'b0;
    wire _112 = 1'b0;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire vdd = 1'b1;
    wire _104 = 1'b0;
    wire _103 = 1'b0;
    wire _102;
    reg _105;
    reg _108;
    reg _111;
    reg _114;
    reg _117;
    reg _120;
    reg _123;
    reg _126;
    reg _129;
    wire _1730;
    wire write_enable_94;
    wire _1735;
    wire gnd = 1'b0;
    wire [131:0] _1742;
    wire [63:0] _1743;
    wire _72;
    wire _1671 = 1'b0;
    wire _1670 = 1'b0;
    wire _1673;
    wire _73;
    reg PHASE_22;
    wire [63:0] _1755;
    wire _76;
    wire _78;
    wire _80;
    wire _82;
    wire _84;
    wire [523:0] _91;
    wire _1756;

    /* logic */
    assign address = _372 ? _199 : _367;
    assign write_enable = _365 & _372;
    assign address_0 = _372 ? _164 : _68;
    assign _374 = ~ _372;
    assign read_enable = _360 & _374;
    assign _372 = ~ PHASE_1;
    assign write_enable_0 = _358 & _372;
    assign _376 = write_enable_0 | read_enable;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_376), .regcea(vdd), .wea(write_enable_0), .addra(address_0), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable), .regceb(vdd), .web(write_enable), .addrb(address), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_381[131:131]), .sbiterrb(_381[130:130]), .doutb(_381[129:66]), .dbiterra(_381[65:65]), .sbiterra(_381[64:64]), .douta(_381[63:0]) );
    assign _382 = _381[63:0];
    assign address_1 = PHASE_1 ? _199 : _367;
    assign _365 = _129 & _328;
    assign write_enable_1 = _365 & PHASE_1;
    assign _279 = _271[129:66];
    assign _278 = _258[129:66];
    assign _280 = PHASE ? _279 : _278;
    assign _276 = _216[129:66];
    assign _275 = _202[129:66];
    assign q1 = PHASE_0 ? _276 : _275;
    assign _281 = _96 ? _280 : q1;
    assign address_2 = _260 ? _254 : _253;
    assign _266 = ~ _260;
    assign read_enable_0 = _102 & _266;
    assign address_3 = _260 ? _60 : _236;
    assign _262 = ~ _260;
    assign read_enable_1 = _102 & _262;
    assign _260 = ~ PHASE;
    assign write_enable_3 = _219 & _260;
    assign _264 = write_enable_3 | read_enable_1;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_0
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_264), .regcea(vdd), .wea(write_enable_3), .addra(address_3), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_0), .regceb(vdd), .web(write_enable_2), .addrb(address_2), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_271[131:131]), .sbiterrb(_271[130:130]), .doutb(_271[129:66]), .dbiterra(_271[65:65]), .sbiterra(_271[64:64]), .douta(_271[63:0]) );
    assign _272 = _271[63:0];
    assign _252 = _172[11:11];
    assign _251 = _172[10:10];
    assign _250 = _172[9:9];
    assign _249 = _172[8:8];
    assign _248 = _172[7:7];
    assign _247 = _172[6:6];
    assign _246 = _172[5:5];
    assign _245 = _172[4:4];
    assign _244 = _172[3:3];
    assign _243 = _172[2:2];
    assign _242 = _172[1:1];
    assign _241 = _172[0:0];
    assign _253 = { _241, _242, _243, _244, _245, _246, _247, _248, _249, _250, _251, _252 };
    assign address_4 = PHASE ? _254 : _253;
    assign _238 = ~ PHASE;
    assign read_enable_2 = _102 & _238;
    assign data_1 = wr_d7;
    assign _235 = _137[11:11];
    assign _234 = _137[10:10];
    assign _233 = _137[9:9];
    assign _232 = _137[8:8];
    assign _231 = _137[7:7];
    assign _230 = _137[6:6];
    assign _229 = _137[5:5];
    assign _228 = _137[4:4];
    assign _227 = _137[3:3];
    assign _226 = _137[2:2];
    assign _225 = _137[1:1];
    assign _224 = _137[0:0];
    assign _236 = { _224, _225, _226, _227, _228, _229, _230, _231, _232, _233, _234, _235 };
    assign address_5 = PHASE ? _60 : _236;
    assign _221 = ~ PHASE;
    assign read_enable_3 = _102 & _221;
    assign _219 = _62[7:7];
    assign write_enable_5 = _219 & PHASE;
    assign _223 = write_enable_5 | read_enable_3;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_1
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_223), .regcea(vdd), .wea(write_enable_5), .addra(address_5), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_2), .regceb(vdd), .web(write_enable_4), .addrb(address_4), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_258[131:131]), .sbiterrb(_258[130:130]), .doutb(_258[129:66]), .dbiterra(_258[65:65]), .sbiterra(_258[64:64]), .douta(_258[63:0]) );
    assign _259 = _258[63:0];
    assign _89 = ~ PHASE;
    assign _3 = _89;
    always @(posedge _84) begin
        if (_82)
            PHASE <= _87;
        else
            if (_72)
                PHASE <= _3;
    end
    assign _273 = PHASE ? _272 : _259;
    assign address_6 = _204 ? _199 : _172;
    assign _211 = ~ _204;
    assign read_enable_4 = _102 & _211;
    assign write_enable_6 = _167 & _204;
    assign _213 = write_enable_6 | read_enable_4;
    assign address_7 = _204 ? _164 : _137;
    assign _206 = ~ _204;
    assign read_enable_5 = _102 & _206;
    assign _204 = ~ PHASE_0;
    assign write_enable_7 = _132 & _204;
    assign _208 = write_enable_7 | read_enable_5;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_2
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_208), .regcea(vdd), .wea(write_enable_7), .addra(address_7), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_213), .regceb(vdd), .web(write_enable_6), .addrb(address_6), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_216[131:131]), .sbiterrb(_216[130:130]), .doutb(_216[129:66]), .dbiterra(_216[65:65]), .sbiterra(_216[64:64]), .douta(_216[63:0]) );
    assign _217 = _216[63:0];
    assign _295 = _294[127:64];
    assign data_3 = _295;
    assign address_8 = PHASE_0 ? _199 : _172;
    assign _169 = ~ PHASE_0;
    assign read_enable_6 = _102 & _169;
    assign _166 = ~ _130;
    assign _167 = _129 & _166;
    assign write_enable_8 = _167 & PHASE_0;
    assign _171 = write_enable_8 | read_enable_6;
    assign address_9 = PHASE_0 ? _164 : _137;
    assign _134 = ~ PHASE_0;
    assign read_enable_7 = _102 & _134;
    assign _131 = ~ _130;
    assign _132 = _129 & _131;
    assign write_enable_9 = _132 & PHASE_0;
    assign _136 = write_enable_9 | read_enable_7;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_3
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_136), .regcea(vdd), .wea(write_enable_9), .addra(address_9), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_171), .regceb(vdd), .web(write_enable_8), .addrb(address_8), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_202[131:131]), .sbiterrb(_202[130:130]), .doutb(_202[129:66]), .dbiterra(_202[65:65]), .sbiterra(_202[64:64]), .douta(_202[63:0]) );
    assign _203 = _202[63:0];
    assign _296 = ~ PHASE_0;
    assign _5 = _296;
    always @(posedge _84) begin
        if (_82)
            PHASE_0 <= _98;
        else
            if (_99)
                PHASE_0 <= _5;
    end
    assign q0 = PHASE_0 ? _217 : _203;
    always @(posedge _84) begin
        if (_82)
            _96 <= _94;
        else
            _96 <= _92;
    end
    assign _274 = _96 ? _273 : q0;
    dp_6
        dp_6
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_274), .d2(_281), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_294[191:128]), .q2(_294[127:64]), .q1(_294[63:0]) );
    assign _297 = _294[63:0];
    assign data_7 = _297;
    assign address_10 = PHASE_1 ? _164 : _68;
    assign _361 = ~ PHASE_1;
    assign _360 = _70[7:7];
    assign read_enable_8 = _360 & _361;
    always @(posedge _84) begin
        if (_82)
            _331 <= _330;
        else
            _331 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _334 <= _333;
        else
            _334 <= _331;
    end
    always @(posedge _84) begin
        if (_82)
            _337 <= _336;
        else
            _337 <= _334;
    end
    always @(posedge _84) begin
        if (_82)
            _340 <= _339;
        else
            _340 <= _337;
    end
    always @(posedge _84) begin
        if (_82)
            _343 <= _342;
        else
            _343 <= _340;
    end
    always @(posedge _84) begin
        if (_82)
            _346 <= _345;
        else
            _346 <= _343;
    end
    always @(posedge _84) begin
        if (_82)
            _349 <= _348;
        else
            _349 <= _346;
    end
    always @(posedge _84) begin
        if (_82)
            _352 <= _351;
        else
            _352 <= _349;
    end
    always @(posedge _84) begin
        if (_82)
            _355 <= _354;
        else
            _355 <= _352;
    end
    assign _356 = ~ _355;
    always @(posedge _84) begin
        if (_82)
            _304 <= _303;
        else
            _304 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _307 <= _306;
        else
            _307 <= _304;
    end
    always @(posedge _84) begin
        if (_82)
            _310 <= _309;
        else
            _310 <= _307;
    end
    always @(posedge _84) begin
        if (_82)
            _313 <= _312;
        else
            _313 <= _310;
    end
    always @(posedge _84) begin
        if (_82)
            _316 <= _315;
        else
            _316 <= _313;
    end
    always @(posedge _84) begin
        if (_82)
            _319 <= _318;
        else
            _319 <= _316;
    end
    always @(posedge _84) begin
        if (_82)
            _322 <= _321;
        else
            _322 <= _319;
    end
    always @(posedge _84) begin
        if (_82)
            _325 <= _324;
        else
            _325 <= _322;
    end
    always @(posedge _84) begin
        if (_82)
            _328 <= _327;
        else
            _328 <= _325;
    end
    assign _357 = _328 & _356;
    assign _358 = _129 & _357;
    assign write_enable_10 = _358 & PHASE_1;
    assign _363 = write_enable_10 | read_enable_8;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_4
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_363), .regcea(vdd), .wea(write_enable_10), .addra(address_10), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_1), .regceb(vdd), .web(write_enable_1), .addrb(address_1), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_370[131:131]), .sbiterrb(_370[130:130]), .doutb(_370[129:66]), .dbiterra(_370[65:65]), .sbiterra(_370[64:64]), .douta(_370[63:0]) );
    assign _371 = _370[63:0];
    assign _301 = ~ PHASE_1;
    assign _7 = _301;
    always @(posedge _84) begin
        if (_82)
            PHASE_1 <= _299;
        else
            if (_72)
                PHASE_1 <= _7;
    end
    assign _383 = PHASE_1 ? _382 : _371;
    assign address_11 = _568 ? _199 : _563;
    assign write_enable_11 = _561 & _568;
    assign address_12 = _568 ? _164 : _68;
    assign _570 = ~ _568;
    assign read_enable_9 = _556 & _570;
    assign _568 = ~ PHASE_4;
    assign write_enable_12 = _554 & _568;
    assign _572 = write_enable_12 | read_enable_9;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_5
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_572), .regcea(vdd), .wea(write_enable_12), .addra(address_12), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_11), .regceb(vdd), .web(write_enable_11), .addrb(address_11), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_577[131:131]), .sbiterrb(_577[130:130]), .doutb(_577[129:66]), .dbiterra(_577[65:65]), .sbiterra(_577[64:64]), .douta(_577[63:0]) );
    assign _578 = _577[63:0];
    assign address_13 = PHASE_4 ? _199 : _563;
    assign _561 = _129 & _524;
    assign write_enable_13 = _561 & PHASE_4;
    assign _486 = _478[129:66];
    assign _485 = _465[129:66];
    assign _487 = PHASE_2 ? _486 : _485;
    assign _483 = _423[129:66];
    assign _482 = _409[129:66];
    assign q1_0 = PHASE_3 ? _483 : _482;
    assign _488 = _390 ? _487 : q1_0;
    assign address_14 = _467 ? _461 : _460;
    assign _473 = ~ _467;
    assign read_enable_10 = _102 & _473;
    assign address_15 = _467 ? _60 : _443;
    assign _469 = ~ _467;
    assign read_enable_11 = _102 & _469;
    assign _467 = ~ PHASE_2;
    assign write_enable_15 = _426 & _467;
    assign _471 = write_enable_15 | read_enable_11;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_6
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_471), .regcea(vdd), .wea(write_enable_15), .addra(address_15), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_10), .regceb(vdd), .web(write_enable_14), .addrb(address_14), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_478[131:131]), .sbiterrb(_478[130:130]), .doutb(_478[129:66]), .dbiterra(_478[65:65]), .sbiterra(_478[64:64]), .douta(_478[63:0]) );
    assign _479 = _478[63:0];
    assign _459 = _172[11:11];
    assign _458 = _172[10:10];
    assign _457 = _172[9:9];
    assign _456 = _172[8:8];
    assign _455 = _172[7:7];
    assign _454 = _172[6:6];
    assign _453 = _172[5:5];
    assign _452 = _172[4:4];
    assign _451 = _172[3:3];
    assign _450 = _172[2:2];
    assign _449 = _172[1:1];
    assign _448 = _172[0:0];
    assign _460 = { _448, _449, _450, _451, _452, _453, _454, _455, _456, _457, _458, _459 };
    assign address_16 = PHASE_2 ? _461 : _460;
    assign _445 = ~ PHASE_2;
    assign read_enable_12 = _102 & _445;
    assign data_13 = wr_d6;
    assign _442 = _137[11:11];
    assign _441 = _137[10:10];
    assign _440 = _137[9:9];
    assign _439 = _137[8:8];
    assign _438 = _137[7:7];
    assign _437 = _137[6:6];
    assign _436 = _137[5:5];
    assign _435 = _137[4:4];
    assign _434 = _137[3:3];
    assign _433 = _137[2:2];
    assign _432 = _137[1:1];
    assign _431 = _137[0:0];
    assign _443 = { _431, _432, _433, _434, _435, _436, _437, _438, _439, _440, _441, _442 };
    assign address_17 = PHASE_2 ? _60 : _443;
    assign _428 = ~ PHASE_2;
    assign read_enable_13 = _102 & _428;
    assign _426 = _62[6:6];
    assign write_enable_17 = _426 & PHASE_2;
    assign _430 = write_enable_17 | read_enable_13;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_7
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_430), .regcea(vdd), .wea(write_enable_17), .addra(address_17), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_12), .regceb(vdd), .web(write_enable_16), .addrb(address_16), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_465[131:131]), .sbiterrb(_465[130:130]), .doutb(_465[129:66]), .dbiterra(_465[65:65]), .sbiterra(_465[64:64]), .douta(_465[63:0]) );
    assign _466 = _465[63:0];
    assign _387 = ~ PHASE_2;
    assign _11 = _387;
    always @(posedge _84) begin
        if (_82)
            PHASE_2 <= _385;
        else
            if (_72)
                PHASE_2 <= _11;
    end
    assign _480 = PHASE_2 ? _479 : _466;
    assign address_18 = _411 ? _199 : _172;
    assign _418 = ~ _411;
    assign read_enable_14 = _102 & _418;
    assign write_enable_18 = _402 & _411;
    assign _420 = write_enable_18 | read_enable_14;
    assign address_19 = _411 ? _164 : _137;
    assign _413 = ~ _411;
    assign read_enable_15 = _102 & _413;
    assign _411 = ~ PHASE_3;
    assign write_enable_19 = _395 & _411;
    assign _415 = write_enable_19 | read_enable_15;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_8
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_415), .regcea(vdd), .wea(write_enable_19), .addra(address_19), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_420), .regceb(vdd), .web(write_enable_18), .addrb(address_18), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_423[131:131]), .sbiterrb(_423[130:130]), .doutb(_423[129:66]), .dbiterra(_423[65:65]), .sbiterra(_423[64:64]), .douta(_423[63:0]) );
    assign _424 = _423[63:0];
    assign _491 = _490[127:64];
    assign data_15 = _491;
    assign address_20 = PHASE_3 ? _199 : _172;
    assign _404 = ~ PHASE_3;
    assign read_enable_16 = _102 & _404;
    assign _401 = ~ _130;
    assign _402 = _129 & _401;
    assign write_enable_20 = _402 & PHASE_3;
    assign _406 = write_enable_20 | read_enable_16;
    assign address_21 = PHASE_3 ? _164 : _137;
    assign _397 = ~ PHASE_3;
    assign read_enable_17 = _102 & _397;
    assign _394 = ~ _130;
    assign _395 = _129 & _394;
    assign write_enable_21 = _395 & PHASE_3;
    assign _399 = write_enable_21 | read_enable_17;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_9
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_399), .regcea(vdd), .wea(write_enable_21), .addra(address_21), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_406), .regceb(vdd), .web(write_enable_20), .addrb(address_20), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_409[131:131]), .sbiterrb(_409[130:130]), .doutb(_409[129:66]), .dbiterra(_409[65:65]), .sbiterra(_409[64:64]), .douta(_409[63:0]) );
    assign _410 = _409[63:0];
    assign _492 = ~ PHASE_3;
    assign _13 = _492;
    always @(posedge _84) begin
        if (_82)
            PHASE_3 <= _392;
        else
            if (_99)
                PHASE_3 <= _13;
    end
    assign q0_0 = PHASE_3 ? _424 : _410;
    always @(posedge _84) begin
        if (_82)
            _390 <= _389;
        else
            _390 <= _92;
    end
    assign _481 = _390 ? _480 : q0_0;
    dp_5
        dp_5
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_481), .d2(_488), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_490[191:128]), .q2(_490[127:64]), .q1(_490[63:0]) );
    assign _493 = _490[63:0];
    assign data_19 = _493;
    assign address_22 = PHASE_4 ? _164 : _68;
    assign _557 = ~ PHASE_4;
    assign _556 = _70[6:6];
    assign read_enable_18 = _556 & _557;
    always @(posedge _84) begin
        if (_82)
            _527 <= _526;
        else
            _527 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _530 <= _529;
        else
            _530 <= _527;
    end
    always @(posedge _84) begin
        if (_82)
            _533 <= _532;
        else
            _533 <= _530;
    end
    always @(posedge _84) begin
        if (_82)
            _536 <= _535;
        else
            _536 <= _533;
    end
    always @(posedge _84) begin
        if (_82)
            _539 <= _538;
        else
            _539 <= _536;
    end
    always @(posedge _84) begin
        if (_82)
            _542 <= _541;
        else
            _542 <= _539;
    end
    always @(posedge _84) begin
        if (_82)
            _545 <= _544;
        else
            _545 <= _542;
    end
    always @(posedge _84) begin
        if (_82)
            _548 <= _547;
        else
            _548 <= _545;
    end
    always @(posedge _84) begin
        if (_82)
            _551 <= _550;
        else
            _551 <= _548;
    end
    assign _552 = ~ _551;
    always @(posedge _84) begin
        if (_82)
            _500 <= _499;
        else
            _500 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _503 <= _502;
        else
            _503 <= _500;
    end
    always @(posedge _84) begin
        if (_82)
            _506 <= _505;
        else
            _506 <= _503;
    end
    always @(posedge _84) begin
        if (_82)
            _509 <= _508;
        else
            _509 <= _506;
    end
    always @(posedge _84) begin
        if (_82)
            _512 <= _511;
        else
            _512 <= _509;
    end
    always @(posedge _84) begin
        if (_82)
            _515 <= _514;
        else
            _515 <= _512;
    end
    always @(posedge _84) begin
        if (_82)
            _518 <= _517;
        else
            _518 <= _515;
    end
    always @(posedge _84) begin
        if (_82)
            _521 <= _520;
        else
            _521 <= _518;
    end
    always @(posedge _84) begin
        if (_82)
            _524 <= _523;
        else
            _524 <= _521;
    end
    assign _553 = _524 & _552;
    assign _554 = _129 & _553;
    assign write_enable_22 = _554 & PHASE_4;
    assign _559 = write_enable_22 | read_enable_18;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_10
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_559), .regcea(vdd), .wea(write_enable_22), .addra(address_22), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_13), .regceb(vdd), .web(write_enable_13), .addrb(address_13), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_566[131:131]), .sbiterrb(_566[130:130]), .doutb(_566[129:66]), .dbiterra(_566[65:65]), .sbiterra(_566[64:64]), .douta(_566[63:0]) );
    assign _567 = _566[63:0];
    assign _497 = ~ PHASE_4;
    assign _15 = _497;
    always @(posedge _84) begin
        if (_82)
            PHASE_4 <= _495;
        else
            if (_72)
                PHASE_4 <= _15;
    end
    assign _579 = PHASE_4 ? _578 : _567;
    assign address_23 = _764 ? _199 : _759;
    assign write_enable_23 = _757 & _764;
    assign address_24 = _764 ? _164 : _68;
    assign _766 = ~ _764;
    assign read_enable_19 = _752 & _766;
    assign _764 = ~ PHASE_7;
    assign write_enable_24 = _750 & _764;
    assign _768 = write_enable_24 | read_enable_19;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_11
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_768), .regcea(vdd), .wea(write_enable_24), .addra(address_24), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_23), .regceb(vdd), .web(write_enable_23), .addrb(address_23), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_773[131:131]), .sbiterrb(_773[130:130]), .doutb(_773[129:66]), .dbiterra(_773[65:65]), .sbiterra(_773[64:64]), .douta(_773[63:0]) );
    assign _774 = _773[63:0];
    assign address_25 = PHASE_7 ? _199 : _759;
    assign _757 = _129 & _720;
    assign write_enable_25 = _757 & PHASE_7;
    assign _682 = _674[129:66];
    assign _681 = _661[129:66];
    assign _683 = PHASE_5 ? _682 : _681;
    assign _679 = _619[129:66];
    assign _678 = _605[129:66];
    assign q1_1 = PHASE_6 ? _679 : _678;
    assign _684 = _586 ? _683 : q1_1;
    assign address_26 = _663 ? _657 : _656;
    assign _669 = ~ _663;
    assign read_enable_20 = _102 & _669;
    assign address_27 = _663 ? _60 : _639;
    assign _665 = ~ _663;
    assign read_enable_21 = _102 & _665;
    assign _663 = ~ PHASE_5;
    assign write_enable_27 = _622 & _663;
    assign _667 = write_enable_27 | read_enable_21;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_12
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_667), .regcea(vdd), .wea(write_enable_27), .addra(address_27), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_20), .regceb(vdd), .web(write_enable_26), .addrb(address_26), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_674[131:131]), .sbiterrb(_674[130:130]), .doutb(_674[129:66]), .dbiterra(_674[65:65]), .sbiterra(_674[64:64]), .douta(_674[63:0]) );
    assign _675 = _674[63:0];
    assign _655 = _172[11:11];
    assign _654 = _172[10:10];
    assign _653 = _172[9:9];
    assign _652 = _172[8:8];
    assign _651 = _172[7:7];
    assign _650 = _172[6:6];
    assign _649 = _172[5:5];
    assign _648 = _172[4:4];
    assign _647 = _172[3:3];
    assign _646 = _172[2:2];
    assign _645 = _172[1:1];
    assign _644 = _172[0:0];
    assign _656 = { _644, _645, _646, _647, _648, _649, _650, _651, _652, _653, _654, _655 };
    assign address_28 = PHASE_5 ? _657 : _656;
    assign _641 = ~ PHASE_5;
    assign read_enable_22 = _102 & _641;
    assign data_25 = wr_d5;
    assign _638 = _137[11:11];
    assign _637 = _137[10:10];
    assign _636 = _137[9:9];
    assign _635 = _137[8:8];
    assign _634 = _137[7:7];
    assign _633 = _137[6:6];
    assign _632 = _137[5:5];
    assign _631 = _137[4:4];
    assign _630 = _137[3:3];
    assign _629 = _137[2:2];
    assign _628 = _137[1:1];
    assign _627 = _137[0:0];
    assign _639 = { _627, _628, _629, _630, _631, _632, _633, _634, _635, _636, _637, _638 };
    assign address_29 = PHASE_5 ? _60 : _639;
    assign _624 = ~ PHASE_5;
    assign read_enable_23 = _102 & _624;
    assign _622 = _62[5:5];
    assign write_enable_29 = _622 & PHASE_5;
    assign _626 = write_enable_29 | read_enable_23;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_13
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_626), .regcea(vdd), .wea(write_enable_29), .addra(address_29), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_22), .regceb(vdd), .web(write_enable_28), .addrb(address_28), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_661[131:131]), .sbiterrb(_661[130:130]), .doutb(_661[129:66]), .dbiterra(_661[65:65]), .sbiterra(_661[64:64]), .douta(_661[63:0]) );
    assign _662 = _661[63:0];
    assign _583 = ~ PHASE_5;
    assign _19 = _583;
    always @(posedge _84) begin
        if (_82)
            PHASE_5 <= _581;
        else
            if (_72)
                PHASE_5 <= _19;
    end
    assign _676 = PHASE_5 ? _675 : _662;
    assign address_30 = _607 ? _199 : _172;
    assign _614 = ~ _607;
    assign read_enable_24 = _102 & _614;
    assign write_enable_30 = _598 & _607;
    assign _616 = write_enable_30 | read_enable_24;
    assign address_31 = _607 ? _164 : _137;
    assign _609 = ~ _607;
    assign read_enable_25 = _102 & _609;
    assign _607 = ~ PHASE_6;
    assign write_enable_31 = _591 & _607;
    assign _611 = write_enable_31 | read_enable_25;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_14
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_611), .regcea(vdd), .wea(write_enable_31), .addra(address_31), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_616), .regceb(vdd), .web(write_enable_30), .addrb(address_30), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_619[131:131]), .sbiterrb(_619[130:130]), .doutb(_619[129:66]), .dbiterra(_619[65:65]), .sbiterra(_619[64:64]), .douta(_619[63:0]) );
    assign _620 = _619[63:0];
    assign _687 = _686[127:64];
    assign data_27 = _687;
    assign address_32 = PHASE_6 ? _199 : _172;
    assign _600 = ~ PHASE_6;
    assign read_enable_26 = _102 & _600;
    assign _597 = ~ _130;
    assign _598 = _129 & _597;
    assign write_enable_32 = _598 & PHASE_6;
    assign _602 = write_enable_32 | read_enable_26;
    assign address_33 = PHASE_6 ? _164 : _137;
    assign _593 = ~ PHASE_6;
    assign read_enable_27 = _102 & _593;
    assign _590 = ~ _130;
    assign _591 = _129 & _590;
    assign write_enable_33 = _591 & PHASE_6;
    assign _595 = write_enable_33 | read_enable_27;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_15
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_595), .regcea(vdd), .wea(write_enable_33), .addra(address_33), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_602), .regceb(vdd), .web(write_enable_32), .addrb(address_32), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_605[131:131]), .sbiterrb(_605[130:130]), .doutb(_605[129:66]), .dbiterra(_605[65:65]), .sbiterra(_605[64:64]), .douta(_605[63:0]) );
    assign _606 = _605[63:0];
    assign _688 = ~ PHASE_6;
    assign _21 = _688;
    always @(posedge _84) begin
        if (_82)
            PHASE_6 <= _588;
        else
            if (_99)
                PHASE_6 <= _21;
    end
    assign q0_1 = PHASE_6 ? _620 : _606;
    always @(posedge _84) begin
        if (_82)
            _586 <= _585;
        else
            _586 <= _92;
    end
    assign _677 = _586 ? _676 : q0_1;
    dp_4
        dp_4
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_677), .d2(_684), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_686[191:128]), .q2(_686[127:64]), .q1(_686[63:0]) );
    assign _689 = _686[63:0];
    assign data_31 = _689;
    assign address_34 = PHASE_7 ? _164 : _68;
    assign _753 = ~ PHASE_7;
    assign _752 = _70[5:5];
    assign read_enable_28 = _752 & _753;
    always @(posedge _84) begin
        if (_82)
            _723 <= _722;
        else
            _723 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _726 <= _725;
        else
            _726 <= _723;
    end
    always @(posedge _84) begin
        if (_82)
            _729 <= _728;
        else
            _729 <= _726;
    end
    always @(posedge _84) begin
        if (_82)
            _732 <= _731;
        else
            _732 <= _729;
    end
    always @(posedge _84) begin
        if (_82)
            _735 <= _734;
        else
            _735 <= _732;
    end
    always @(posedge _84) begin
        if (_82)
            _738 <= _737;
        else
            _738 <= _735;
    end
    always @(posedge _84) begin
        if (_82)
            _741 <= _740;
        else
            _741 <= _738;
    end
    always @(posedge _84) begin
        if (_82)
            _744 <= _743;
        else
            _744 <= _741;
    end
    always @(posedge _84) begin
        if (_82)
            _747 <= _746;
        else
            _747 <= _744;
    end
    assign _748 = ~ _747;
    always @(posedge _84) begin
        if (_82)
            _696 <= _695;
        else
            _696 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _699 <= _698;
        else
            _699 <= _696;
    end
    always @(posedge _84) begin
        if (_82)
            _702 <= _701;
        else
            _702 <= _699;
    end
    always @(posedge _84) begin
        if (_82)
            _705 <= _704;
        else
            _705 <= _702;
    end
    always @(posedge _84) begin
        if (_82)
            _708 <= _707;
        else
            _708 <= _705;
    end
    always @(posedge _84) begin
        if (_82)
            _711 <= _710;
        else
            _711 <= _708;
    end
    always @(posedge _84) begin
        if (_82)
            _714 <= _713;
        else
            _714 <= _711;
    end
    always @(posedge _84) begin
        if (_82)
            _717 <= _716;
        else
            _717 <= _714;
    end
    always @(posedge _84) begin
        if (_82)
            _720 <= _719;
        else
            _720 <= _717;
    end
    assign _749 = _720 & _748;
    assign _750 = _129 & _749;
    assign write_enable_34 = _750 & PHASE_7;
    assign _755 = write_enable_34 | read_enable_28;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_16
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_755), .regcea(vdd), .wea(write_enable_34), .addra(address_34), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_25), .regceb(vdd), .web(write_enable_25), .addrb(address_25), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_762[131:131]), .sbiterrb(_762[130:130]), .doutb(_762[129:66]), .dbiterra(_762[65:65]), .sbiterra(_762[64:64]), .douta(_762[63:0]) );
    assign _763 = _762[63:0];
    assign _693 = ~ PHASE_7;
    assign _23 = _693;
    always @(posedge _84) begin
        if (_82)
            PHASE_7 <= _691;
        else
            if (_72)
                PHASE_7 <= _23;
    end
    assign _775 = PHASE_7 ? _774 : _763;
    assign address_35 = _960 ? _199 : _955;
    assign write_enable_35 = _953 & _960;
    assign address_36 = _960 ? _164 : _68;
    assign _962 = ~ _960;
    assign read_enable_29 = _948 & _962;
    assign _960 = ~ PHASE_10;
    assign write_enable_36 = _946 & _960;
    assign _964 = write_enable_36 | read_enable_29;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_17
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_964), .regcea(vdd), .wea(write_enable_36), .addra(address_36), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_35), .regceb(vdd), .web(write_enable_35), .addrb(address_35), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_969[131:131]), .sbiterrb(_969[130:130]), .doutb(_969[129:66]), .dbiterra(_969[65:65]), .sbiterra(_969[64:64]), .douta(_969[63:0]) );
    assign _970 = _969[63:0];
    assign address_37 = PHASE_10 ? _199 : _955;
    assign _953 = _129 & _916;
    assign write_enable_37 = _953 & PHASE_10;
    assign _878 = _870[129:66];
    assign _877 = _857[129:66];
    assign _879 = PHASE_8 ? _878 : _877;
    assign _875 = _815[129:66];
    assign _874 = _801[129:66];
    assign q1_2 = PHASE_9 ? _875 : _874;
    assign _880 = _782 ? _879 : q1_2;
    assign address_38 = _859 ? _853 : _852;
    assign _865 = ~ _859;
    assign read_enable_30 = _102 & _865;
    assign address_39 = _859 ? _60 : _835;
    assign _861 = ~ _859;
    assign read_enable_31 = _102 & _861;
    assign _859 = ~ PHASE_8;
    assign write_enable_39 = _818 & _859;
    assign _863 = write_enable_39 | read_enable_31;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_18
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_863), .regcea(vdd), .wea(write_enable_39), .addra(address_39), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_30), .regceb(vdd), .web(write_enable_38), .addrb(address_38), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_870[131:131]), .sbiterrb(_870[130:130]), .doutb(_870[129:66]), .dbiterra(_870[65:65]), .sbiterra(_870[64:64]), .douta(_870[63:0]) );
    assign _871 = _870[63:0];
    assign _851 = _172[11:11];
    assign _850 = _172[10:10];
    assign _849 = _172[9:9];
    assign _848 = _172[8:8];
    assign _847 = _172[7:7];
    assign _846 = _172[6:6];
    assign _845 = _172[5:5];
    assign _844 = _172[4:4];
    assign _843 = _172[3:3];
    assign _842 = _172[2:2];
    assign _841 = _172[1:1];
    assign _840 = _172[0:0];
    assign _852 = { _840, _841, _842, _843, _844, _845, _846, _847, _848, _849, _850, _851 };
    assign address_40 = PHASE_8 ? _853 : _852;
    assign _837 = ~ PHASE_8;
    assign read_enable_32 = _102 & _837;
    assign data_37 = wr_d4;
    assign _834 = _137[11:11];
    assign _833 = _137[10:10];
    assign _832 = _137[9:9];
    assign _831 = _137[8:8];
    assign _830 = _137[7:7];
    assign _829 = _137[6:6];
    assign _828 = _137[5:5];
    assign _827 = _137[4:4];
    assign _826 = _137[3:3];
    assign _825 = _137[2:2];
    assign _824 = _137[1:1];
    assign _823 = _137[0:0];
    assign _835 = { _823, _824, _825, _826, _827, _828, _829, _830, _831, _832, _833, _834 };
    assign address_41 = PHASE_8 ? _60 : _835;
    assign _820 = ~ PHASE_8;
    assign read_enable_33 = _102 & _820;
    assign _818 = _62[4:4];
    assign write_enable_41 = _818 & PHASE_8;
    assign _822 = write_enable_41 | read_enable_33;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_19
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_822), .regcea(vdd), .wea(write_enable_41), .addra(address_41), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_32), .regceb(vdd), .web(write_enable_40), .addrb(address_40), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_857[131:131]), .sbiterrb(_857[130:130]), .doutb(_857[129:66]), .dbiterra(_857[65:65]), .sbiterra(_857[64:64]), .douta(_857[63:0]) );
    assign _858 = _857[63:0];
    assign _779 = ~ PHASE_8;
    assign _27 = _779;
    always @(posedge _84) begin
        if (_82)
            PHASE_8 <= _777;
        else
            if (_72)
                PHASE_8 <= _27;
    end
    assign _872 = PHASE_8 ? _871 : _858;
    assign address_42 = _803 ? _199 : _172;
    assign _810 = ~ _803;
    assign read_enable_34 = _102 & _810;
    assign write_enable_42 = _794 & _803;
    assign _812 = write_enable_42 | read_enable_34;
    assign address_43 = _803 ? _164 : _137;
    assign _805 = ~ _803;
    assign read_enable_35 = _102 & _805;
    assign _803 = ~ PHASE_9;
    assign write_enable_43 = _787 & _803;
    assign _807 = write_enable_43 | read_enable_35;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_20
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_807), .regcea(vdd), .wea(write_enable_43), .addra(address_43), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_812), .regceb(vdd), .web(write_enable_42), .addrb(address_42), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_815[131:131]), .sbiterrb(_815[130:130]), .doutb(_815[129:66]), .dbiterra(_815[65:65]), .sbiterra(_815[64:64]), .douta(_815[63:0]) );
    assign _816 = _815[63:0];
    assign _883 = _882[127:64];
    assign data_39 = _883;
    assign address_44 = PHASE_9 ? _199 : _172;
    assign _796 = ~ PHASE_9;
    assign read_enable_36 = _102 & _796;
    assign _793 = ~ _130;
    assign _794 = _129 & _793;
    assign write_enable_44 = _794 & PHASE_9;
    assign _798 = write_enable_44 | read_enable_36;
    assign address_45 = PHASE_9 ? _164 : _137;
    assign _789 = ~ PHASE_9;
    assign read_enable_37 = _102 & _789;
    assign _786 = ~ _130;
    assign _787 = _129 & _786;
    assign write_enable_45 = _787 & PHASE_9;
    assign _791 = write_enable_45 | read_enable_37;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_21
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_791), .regcea(vdd), .wea(write_enable_45), .addra(address_45), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_798), .regceb(vdd), .web(write_enable_44), .addrb(address_44), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_801[131:131]), .sbiterrb(_801[130:130]), .doutb(_801[129:66]), .dbiterra(_801[65:65]), .sbiterra(_801[64:64]), .douta(_801[63:0]) );
    assign _802 = _801[63:0];
    assign _884 = ~ PHASE_9;
    assign _29 = _884;
    always @(posedge _84) begin
        if (_82)
            PHASE_9 <= _784;
        else
            if (_99)
                PHASE_9 <= _29;
    end
    assign q0_2 = PHASE_9 ? _816 : _802;
    always @(posedge _84) begin
        if (_82)
            _782 <= _781;
        else
            _782 <= _92;
    end
    assign _873 = _782 ? _872 : q0_2;
    dp_3
        dp_3
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_873), .d2(_880), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_882[191:128]), .q2(_882[127:64]), .q1(_882[63:0]) );
    assign _885 = _882[63:0];
    assign data_43 = _885;
    assign address_46 = PHASE_10 ? _164 : _68;
    assign _949 = ~ PHASE_10;
    assign _948 = _70[4:4];
    assign read_enable_38 = _948 & _949;
    always @(posedge _84) begin
        if (_82)
            _919 <= _918;
        else
            _919 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _922 <= _921;
        else
            _922 <= _919;
    end
    always @(posedge _84) begin
        if (_82)
            _925 <= _924;
        else
            _925 <= _922;
    end
    always @(posedge _84) begin
        if (_82)
            _928 <= _927;
        else
            _928 <= _925;
    end
    always @(posedge _84) begin
        if (_82)
            _931 <= _930;
        else
            _931 <= _928;
    end
    always @(posedge _84) begin
        if (_82)
            _934 <= _933;
        else
            _934 <= _931;
    end
    always @(posedge _84) begin
        if (_82)
            _937 <= _936;
        else
            _937 <= _934;
    end
    always @(posedge _84) begin
        if (_82)
            _940 <= _939;
        else
            _940 <= _937;
    end
    always @(posedge _84) begin
        if (_82)
            _943 <= _942;
        else
            _943 <= _940;
    end
    assign _944 = ~ _943;
    always @(posedge _84) begin
        if (_82)
            _892 <= _891;
        else
            _892 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _895 <= _894;
        else
            _895 <= _892;
    end
    always @(posedge _84) begin
        if (_82)
            _898 <= _897;
        else
            _898 <= _895;
    end
    always @(posedge _84) begin
        if (_82)
            _901 <= _900;
        else
            _901 <= _898;
    end
    always @(posedge _84) begin
        if (_82)
            _904 <= _903;
        else
            _904 <= _901;
    end
    always @(posedge _84) begin
        if (_82)
            _907 <= _906;
        else
            _907 <= _904;
    end
    always @(posedge _84) begin
        if (_82)
            _910 <= _909;
        else
            _910 <= _907;
    end
    always @(posedge _84) begin
        if (_82)
            _913 <= _912;
        else
            _913 <= _910;
    end
    always @(posedge _84) begin
        if (_82)
            _916 <= _915;
        else
            _916 <= _913;
    end
    assign _945 = _916 & _944;
    assign _946 = _129 & _945;
    assign write_enable_46 = _946 & PHASE_10;
    assign _951 = write_enable_46 | read_enable_38;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_22
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_951), .regcea(vdd), .wea(write_enable_46), .addra(address_46), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_37), .regceb(vdd), .web(write_enable_37), .addrb(address_37), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_958[131:131]), .sbiterrb(_958[130:130]), .doutb(_958[129:66]), .dbiterra(_958[65:65]), .sbiterra(_958[64:64]), .douta(_958[63:0]) );
    assign _959 = _958[63:0];
    assign _889 = ~ PHASE_10;
    assign _31 = _889;
    always @(posedge _84) begin
        if (_82)
            PHASE_10 <= _887;
        else
            if (_72)
                PHASE_10 <= _31;
    end
    assign _971 = PHASE_10 ? _970 : _959;
    assign address_47 = _1156 ? _199 : _1151;
    assign write_enable_47 = _1149 & _1156;
    assign address_48 = _1156 ? _164 : _68;
    assign _1158 = ~ _1156;
    assign read_enable_39 = _1144 & _1158;
    assign _1156 = ~ PHASE_13;
    assign write_enable_48 = _1142 & _1156;
    assign _1160 = write_enable_48 | read_enable_39;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_23
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1160), .regcea(vdd), .wea(write_enable_48), .addra(address_48), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_47), .regceb(vdd), .web(write_enable_47), .addrb(address_47), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1165[131:131]), .sbiterrb(_1165[130:130]), .doutb(_1165[129:66]), .dbiterra(_1165[65:65]), .sbiterra(_1165[64:64]), .douta(_1165[63:0]) );
    assign _1166 = _1165[63:0];
    assign address_49 = PHASE_13 ? _199 : _1151;
    assign _1149 = _129 & _1112;
    assign write_enable_49 = _1149 & PHASE_13;
    assign _1074 = _1066[129:66];
    assign _1073 = _1053[129:66];
    assign _1075 = PHASE_11 ? _1074 : _1073;
    assign _1071 = _1011[129:66];
    assign _1070 = _997[129:66];
    assign q1_3 = PHASE_12 ? _1071 : _1070;
    assign _1076 = _978 ? _1075 : q1_3;
    assign address_50 = _1055 ? _1049 : _1048;
    assign _1061 = ~ _1055;
    assign read_enable_40 = _102 & _1061;
    assign address_51 = _1055 ? _60 : _1031;
    assign _1057 = ~ _1055;
    assign read_enable_41 = _102 & _1057;
    assign _1055 = ~ PHASE_11;
    assign write_enable_51 = _1014 & _1055;
    assign _1059 = write_enable_51 | read_enable_41;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_24
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1059), .regcea(vdd), .wea(write_enable_51), .addra(address_51), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_40), .regceb(vdd), .web(write_enable_50), .addrb(address_50), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1066[131:131]), .sbiterrb(_1066[130:130]), .doutb(_1066[129:66]), .dbiterra(_1066[65:65]), .sbiterra(_1066[64:64]), .douta(_1066[63:0]) );
    assign _1067 = _1066[63:0];
    assign _1047 = _172[11:11];
    assign _1046 = _172[10:10];
    assign _1045 = _172[9:9];
    assign _1044 = _172[8:8];
    assign _1043 = _172[7:7];
    assign _1042 = _172[6:6];
    assign _1041 = _172[5:5];
    assign _1040 = _172[4:4];
    assign _1039 = _172[3:3];
    assign _1038 = _172[2:2];
    assign _1037 = _172[1:1];
    assign _1036 = _172[0:0];
    assign _1048 = { _1036, _1037, _1038, _1039, _1040, _1041, _1042, _1043, _1044, _1045, _1046, _1047 };
    assign address_52 = PHASE_11 ? _1049 : _1048;
    assign _1033 = ~ PHASE_11;
    assign read_enable_42 = _102 & _1033;
    assign data_49 = wr_d3;
    assign _1030 = _137[11:11];
    assign _1029 = _137[10:10];
    assign _1028 = _137[9:9];
    assign _1027 = _137[8:8];
    assign _1026 = _137[7:7];
    assign _1025 = _137[6:6];
    assign _1024 = _137[5:5];
    assign _1023 = _137[4:4];
    assign _1022 = _137[3:3];
    assign _1021 = _137[2:2];
    assign _1020 = _137[1:1];
    assign _1019 = _137[0:0];
    assign _1031 = { _1019, _1020, _1021, _1022, _1023, _1024, _1025, _1026, _1027, _1028, _1029, _1030 };
    assign address_53 = PHASE_11 ? _60 : _1031;
    assign _1016 = ~ PHASE_11;
    assign read_enable_43 = _102 & _1016;
    assign _1014 = _62[3:3];
    assign write_enable_53 = _1014 & PHASE_11;
    assign _1018 = write_enable_53 | read_enable_43;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_25
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1018), .regcea(vdd), .wea(write_enable_53), .addra(address_53), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_42), .regceb(vdd), .web(write_enable_52), .addrb(address_52), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1053[131:131]), .sbiterrb(_1053[130:130]), .doutb(_1053[129:66]), .dbiterra(_1053[65:65]), .sbiterra(_1053[64:64]), .douta(_1053[63:0]) );
    assign _1054 = _1053[63:0];
    assign _975 = ~ PHASE_11;
    assign _35 = _975;
    always @(posedge _84) begin
        if (_82)
            PHASE_11 <= _973;
        else
            if (_72)
                PHASE_11 <= _35;
    end
    assign _1068 = PHASE_11 ? _1067 : _1054;
    assign address_54 = _999 ? _199 : _172;
    assign _1006 = ~ _999;
    assign read_enable_44 = _102 & _1006;
    assign write_enable_54 = _990 & _999;
    assign _1008 = write_enable_54 | read_enable_44;
    assign address_55 = _999 ? _164 : _137;
    assign _1001 = ~ _999;
    assign read_enable_45 = _102 & _1001;
    assign _999 = ~ PHASE_12;
    assign write_enable_55 = _983 & _999;
    assign _1003 = write_enable_55 | read_enable_45;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_26
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1003), .regcea(vdd), .wea(write_enable_55), .addra(address_55), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1008), .regceb(vdd), .web(write_enable_54), .addrb(address_54), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1011[131:131]), .sbiterrb(_1011[130:130]), .doutb(_1011[129:66]), .dbiterra(_1011[65:65]), .sbiterra(_1011[64:64]), .douta(_1011[63:0]) );
    assign _1012 = _1011[63:0];
    assign _1079 = _1078[127:64];
    assign data_51 = _1079;
    assign address_56 = PHASE_12 ? _199 : _172;
    assign _992 = ~ PHASE_12;
    assign read_enable_46 = _102 & _992;
    assign _989 = ~ _130;
    assign _990 = _129 & _989;
    assign write_enable_56 = _990 & PHASE_12;
    assign _994 = write_enable_56 | read_enable_46;
    assign address_57 = PHASE_12 ? _164 : _137;
    assign _985 = ~ PHASE_12;
    assign read_enable_47 = _102 & _985;
    assign _982 = ~ _130;
    assign _983 = _129 & _982;
    assign write_enable_57 = _983 & PHASE_12;
    assign _987 = write_enable_57 | read_enable_47;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_27
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_987), .regcea(vdd), .wea(write_enable_57), .addra(address_57), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_994), .regceb(vdd), .web(write_enable_56), .addrb(address_56), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_997[131:131]), .sbiterrb(_997[130:130]), .doutb(_997[129:66]), .dbiterra(_997[65:65]), .sbiterra(_997[64:64]), .douta(_997[63:0]) );
    assign _998 = _997[63:0];
    assign _1080 = ~ PHASE_12;
    assign _37 = _1080;
    always @(posedge _84) begin
        if (_82)
            PHASE_12 <= _980;
        else
            if (_99)
                PHASE_12 <= _37;
    end
    assign q0_3 = PHASE_12 ? _1012 : _998;
    always @(posedge _84) begin
        if (_82)
            _978 <= _977;
        else
            _978 <= _92;
    end
    assign _1069 = _978 ? _1068 : q0_3;
    dp_2
        dp_2
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1069), .d2(_1076), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1078[191:128]), .q2(_1078[127:64]), .q1(_1078[63:0]) );
    assign _1081 = _1078[63:0];
    assign data_55 = _1081;
    assign address_58 = PHASE_13 ? _164 : _68;
    assign _1145 = ~ PHASE_13;
    assign _1144 = _70[3:3];
    assign read_enable_48 = _1144 & _1145;
    always @(posedge _84) begin
        if (_82)
            _1115 <= _1114;
        else
            _1115 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1118 <= _1117;
        else
            _1118 <= _1115;
    end
    always @(posedge _84) begin
        if (_82)
            _1121 <= _1120;
        else
            _1121 <= _1118;
    end
    always @(posedge _84) begin
        if (_82)
            _1124 <= _1123;
        else
            _1124 <= _1121;
    end
    always @(posedge _84) begin
        if (_82)
            _1127 <= _1126;
        else
            _1127 <= _1124;
    end
    always @(posedge _84) begin
        if (_82)
            _1130 <= _1129;
        else
            _1130 <= _1127;
    end
    always @(posedge _84) begin
        if (_82)
            _1133 <= _1132;
        else
            _1133 <= _1130;
    end
    always @(posedge _84) begin
        if (_82)
            _1136 <= _1135;
        else
            _1136 <= _1133;
    end
    always @(posedge _84) begin
        if (_82)
            _1139 <= _1138;
        else
            _1139 <= _1136;
    end
    assign _1140 = ~ _1139;
    always @(posedge _84) begin
        if (_82)
            _1088 <= _1087;
        else
            _1088 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1091 <= _1090;
        else
            _1091 <= _1088;
    end
    always @(posedge _84) begin
        if (_82)
            _1094 <= _1093;
        else
            _1094 <= _1091;
    end
    always @(posedge _84) begin
        if (_82)
            _1097 <= _1096;
        else
            _1097 <= _1094;
    end
    always @(posedge _84) begin
        if (_82)
            _1100 <= _1099;
        else
            _1100 <= _1097;
    end
    always @(posedge _84) begin
        if (_82)
            _1103 <= _1102;
        else
            _1103 <= _1100;
    end
    always @(posedge _84) begin
        if (_82)
            _1106 <= _1105;
        else
            _1106 <= _1103;
    end
    always @(posedge _84) begin
        if (_82)
            _1109 <= _1108;
        else
            _1109 <= _1106;
    end
    always @(posedge _84) begin
        if (_82)
            _1112 <= _1111;
        else
            _1112 <= _1109;
    end
    assign _1141 = _1112 & _1140;
    assign _1142 = _129 & _1141;
    assign write_enable_58 = _1142 & PHASE_13;
    assign _1147 = write_enable_58 | read_enable_48;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_28
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1147), .regcea(vdd), .wea(write_enable_58), .addra(address_58), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_49), .regceb(vdd), .web(write_enable_49), .addrb(address_49), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1154[131:131]), .sbiterrb(_1154[130:130]), .doutb(_1154[129:66]), .dbiterra(_1154[65:65]), .sbiterra(_1154[64:64]), .douta(_1154[63:0]) );
    assign _1155 = _1154[63:0];
    assign _1085 = ~ PHASE_13;
    assign _39 = _1085;
    always @(posedge _84) begin
        if (_82)
            PHASE_13 <= _1083;
        else
            if (_72)
                PHASE_13 <= _39;
    end
    assign _1167 = PHASE_13 ? _1166 : _1155;
    assign address_59 = _1352 ? _199 : _1347;
    assign write_enable_59 = _1345 & _1352;
    assign address_60 = _1352 ? _164 : _68;
    assign _1354 = ~ _1352;
    assign read_enable_49 = _1340 & _1354;
    assign _1352 = ~ PHASE_16;
    assign write_enable_60 = _1338 & _1352;
    assign _1356 = write_enable_60 | read_enable_49;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_29
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1356), .regcea(vdd), .wea(write_enable_60), .addra(address_60), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_59), .regceb(vdd), .web(write_enable_59), .addrb(address_59), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1361[131:131]), .sbiterrb(_1361[130:130]), .doutb(_1361[129:66]), .dbiterra(_1361[65:65]), .sbiterra(_1361[64:64]), .douta(_1361[63:0]) );
    assign _1362 = _1361[63:0];
    assign address_61 = PHASE_16 ? _199 : _1347;
    assign _1345 = _129 & _1308;
    assign write_enable_61 = _1345 & PHASE_16;
    assign _1270 = _1262[129:66];
    assign _1269 = _1249[129:66];
    assign _1271 = PHASE_14 ? _1270 : _1269;
    assign _1267 = _1207[129:66];
    assign _1266 = _1193[129:66];
    assign q1_4 = PHASE_15 ? _1267 : _1266;
    assign _1272 = _1174 ? _1271 : q1_4;
    assign address_62 = _1251 ? _1245 : _1244;
    assign _1257 = ~ _1251;
    assign read_enable_50 = _102 & _1257;
    assign address_63 = _1251 ? _60 : _1227;
    assign _1253 = ~ _1251;
    assign read_enable_51 = _102 & _1253;
    assign _1251 = ~ PHASE_14;
    assign write_enable_63 = _1210 & _1251;
    assign _1255 = write_enable_63 | read_enable_51;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_30
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1255), .regcea(vdd), .wea(write_enable_63), .addra(address_63), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_50), .regceb(vdd), .web(write_enable_62), .addrb(address_62), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1262[131:131]), .sbiterrb(_1262[130:130]), .doutb(_1262[129:66]), .dbiterra(_1262[65:65]), .sbiterra(_1262[64:64]), .douta(_1262[63:0]) );
    assign _1263 = _1262[63:0];
    assign _1243 = _172[11:11];
    assign _1242 = _172[10:10];
    assign _1241 = _172[9:9];
    assign _1240 = _172[8:8];
    assign _1239 = _172[7:7];
    assign _1238 = _172[6:6];
    assign _1237 = _172[5:5];
    assign _1236 = _172[4:4];
    assign _1235 = _172[3:3];
    assign _1234 = _172[2:2];
    assign _1233 = _172[1:1];
    assign _1232 = _172[0:0];
    assign _1244 = { _1232, _1233, _1234, _1235, _1236, _1237, _1238, _1239, _1240, _1241, _1242, _1243 };
    assign address_64 = PHASE_14 ? _1245 : _1244;
    assign _1229 = ~ PHASE_14;
    assign read_enable_52 = _102 & _1229;
    assign data_61 = wr_d2;
    assign _1226 = _137[11:11];
    assign _1225 = _137[10:10];
    assign _1224 = _137[9:9];
    assign _1223 = _137[8:8];
    assign _1222 = _137[7:7];
    assign _1221 = _137[6:6];
    assign _1220 = _137[5:5];
    assign _1219 = _137[4:4];
    assign _1218 = _137[3:3];
    assign _1217 = _137[2:2];
    assign _1216 = _137[1:1];
    assign _1215 = _137[0:0];
    assign _1227 = { _1215, _1216, _1217, _1218, _1219, _1220, _1221, _1222, _1223, _1224, _1225, _1226 };
    assign address_65 = PHASE_14 ? _60 : _1227;
    assign _1212 = ~ PHASE_14;
    assign read_enable_53 = _102 & _1212;
    assign _1210 = _62[2:2];
    assign write_enable_65 = _1210 & PHASE_14;
    assign _1214 = write_enable_65 | read_enable_53;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_31
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1214), .regcea(vdd), .wea(write_enable_65), .addra(address_65), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_52), .regceb(vdd), .web(write_enable_64), .addrb(address_64), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1249[131:131]), .sbiterrb(_1249[130:130]), .doutb(_1249[129:66]), .dbiterra(_1249[65:65]), .sbiterra(_1249[64:64]), .douta(_1249[63:0]) );
    assign _1250 = _1249[63:0];
    assign _1171 = ~ PHASE_14;
    assign _43 = _1171;
    always @(posedge _84) begin
        if (_82)
            PHASE_14 <= _1169;
        else
            if (_72)
                PHASE_14 <= _43;
    end
    assign _1264 = PHASE_14 ? _1263 : _1250;
    assign address_66 = _1195 ? _199 : _172;
    assign _1202 = ~ _1195;
    assign read_enable_54 = _102 & _1202;
    assign write_enable_66 = _1186 & _1195;
    assign _1204 = write_enable_66 | read_enable_54;
    assign address_67 = _1195 ? _164 : _137;
    assign _1197 = ~ _1195;
    assign read_enable_55 = _102 & _1197;
    assign _1195 = ~ PHASE_15;
    assign write_enable_67 = _1179 & _1195;
    assign _1199 = write_enable_67 | read_enable_55;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_32
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1199), .regcea(vdd), .wea(write_enable_67), .addra(address_67), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1204), .regceb(vdd), .web(write_enable_66), .addrb(address_66), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1207[131:131]), .sbiterrb(_1207[130:130]), .doutb(_1207[129:66]), .dbiterra(_1207[65:65]), .sbiterra(_1207[64:64]), .douta(_1207[63:0]) );
    assign _1208 = _1207[63:0];
    assign _1275 = _1274[127:64];
    assign data_63 = _1275;
    assign address_68 = PHASE_15 ? _199 : _172;
    assign _1188 = ~ PHASE_15;
    assign read_enable_56 = _102 & _1188;
    assign _1185 = ~ _130;
    assign _1186 = _129 & _1185;
    assign write_enable_68 = _1186 & PHASE_15;
    assign _1190 = write_enable_68 | read_enable_56;
    assign address_69 = PHASE_15 ? _164 : _137;
    assign _1181 = ~ PHASE_15;
    assign read_enable_57 = _102 & _1181;
    assign _1178 = ~ _130;
    assign _1179 = _129 & _1178;
    assign write_enable_69 = _1179 & PHASE_15;
    assign _1183 = write_enable_69 | read_enable_57;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_33
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1183), .regcea(vdd), .wea(write_enable_69), .addra(address_69), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1190), .regceb(vdd), .web(write_enable_68), .addrb(address_68), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1193[131:131]), .sbiterrb(_1193[130:130]), .doutb(_1193[129:66]), .dbiterra(_1193[65:65]), .sbiterra(_1193[64:64]), .douta(_1193[63:0]) );
    assign _1194 = _1193[63:0];
    assign _1276 = ~ PHASE_15;
    assign _45 = _1276;
    always @(posedge _84) begin
        if (_82)
            PHASE_15 <= _1176;
        else
            if (_99)
                PHASE_15 <= _45;
    end
    assign q0_4 = PHASE_15 ? _1208 : _1194;
    always @(posedge _84) begin
        if (_82)
            _1174 <= _1173;
        else
            _1174 <= _92;
    end
    assign _1265 = _1174 ? _1264 : q0_4;
    dp_1
        dp_1
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1265), .d2(_1272), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1274[191:128]), .q2(_1274[127:64]), .q1(_1274[63:0]) );
    assign _1277 = _1274[63:0];
    assign data_67 = _1277;
    assign address_70 = PHASE_16 ? _164 : _68;
    assign _1341 = ~ PHASE_16;
    assign _1340 = _70[2:2];
    assign read_enable_58 = _1340 & _1341;
    always @(posedge _84) begin
        if (_82)
            _1311 <= _1310;
        else
            _1311 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1314 <= _1313;
        else
            _1314 <= _1311;
    end
    always @(posedge _84) begin
        if (_82)
            _1317 <= _1316;
        else
            _1317 <= _1314;
    end
    always @(posedge _84) begin
        if (_82)
            _1320 <= _1319;
        else
            _1320 <= _1317;
    end
    always @(posedge _84) begin
        if (_82)
            _1323 <= _1322;
        else
            _1323 <= _1320;
    end
    always @(posedge _84) begin
        if (_82)
            _1326 <= _1325;
        else
            _1326 <= _1323;
    end
    always @(posedge _84) begin
        if (_82)
            _1329 <= _1328;
        else
            _1329 <= _1326;
    end
    always @(posedge _84) begin
        if (_82)
            _1332 <= _1331;
        else
            _1332 <= _1329;
    end
    always @(posedge _84) begin
        if (_82)
            _1335 <= _1334;
        else
            _1335 <= _1332;
    end
    assign _1336 = ~ _1335;
    always @(posedge _84) begin
        if (_82)
            _1284 <= _1283;
        else
            _1284 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1287 <= _1286;
        else
            _1287 <= _1284;
    end
    always @(posedge _84) begin
        if (_82)
            _1290 <= _1289;
        else
            _1290 <= _1287;
    end
    always @(posedge _84) begin
        if (_82)
            _1293 <= _1292;
        else
            _1293 <= _1290;
    end
    always @(posedge _84) begin
        if (_82)
            _1296 <= _1295;
        else
            _1296 <= _1293;
    end
    always @(posedge _84) begin
        if (_82)
            _1299 <= _1298;
        else
            _1299 <= _1296;
    end
    always @(posedge _84) begin
        if (_82)
            _1302 <= _1301;
        else
            _1302 <= _1299;
    end
    always @(posedge _84) begin
        if (_82)
            _1305 <= _1304;
        else
            _1305 <= _1302;
    end
    always @(posedge _84) begin
        if (_82)
            _1308 <= _1307;
        else
            _1308 <= _1305;
    end
    assign _1337 = _1308 & _1336;
    assign _1338 = _129 & _1337;
    assign write_enable_70 = _1338 & PHASE_16;
    assign _1343 = write_enable_70 | read_enable_58;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_34
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1343), .regcea(vdd), .wea(write_enable_70), .addra(address_70), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_61), .regceb(vdd), .web(write_enable_61), .addrb(address_61), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1350[131:131]), .sbiterrb(_1350[130:130]), .doutb(_1350[129:66]), .dbiterra(_1350[65:65]), .sbiterra(_1350[64:64]), .douta(_1350[63:0]) );
    assign _1351 = _1350[63:0];
    assign _1281 = ~ PHASE_16;
    assign _47 = _1281;
    always @(posedge _84) begin
        if (_82)
            PHASE_16 <= _1279;
        else
            if (_72)
                PHASE_16 <= _47;
    end
    assign _1363 = PHASE_16 ? _1362 : _1351;
    assign address_71 = _1548 ? _199 : _1543;
    assign write_enable_71 = _1541 & _1548;
    assign address_72 = _1548 ? _164 : _68;
    assign _1550 = ~ _1548;
    assign read_enable_59 = _1536 & _1550;
    assign _1548 = ~ PHASE_19;
    assign write_enable_72 = _1534 & _1548;
    assign _1552 = write_enable_72 | read_enable_59;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_35
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1552), .regcea(vdd), .wea(write_enable_72), .addra(address_72), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_71), .regceb(vdd), .web(write_enable_71), .addrb(address_71), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1557[131:131]), .sbiterrb(_1557[130:130]), .doutb(_1557[129:66]), .dbiterra(_1557[65:65]), .sbiterra(_1557[64:64]), .douta(_1557[63:0]) );
    assign _1558 = _1557[63:0];
    assign address_73 = PHASE_19 ? _199 : _1543;
    assign _1541 = _129 & _1504;
    assign write_enable_73 = _1541 & PHASE_19;
    assign _1466 = _1458[129:66];
    assign _1465 = _1445[129:66];
    assign _1467 = PHASE_17 ? _1466 : _1465;
    assign _1463 = _1403[129:66];
    assign _1462 = _1389[129:66];
    assign q1_5 = PHASE_18 ? _1463 : _1462;
    assign _1468 = _1370 ? _1467 : q1_5;
    assign address_74 = _1447 ? _1441 : _1440;
    assign _1453 = ~ _1447;
    assign read_enable_60 = _102 & _1453;
    assign address_75 = _1447 ? _60 : _1423;
    assign _1449 = ~ _1447;
    assign read_enable_61 = _102 & _1449;
    assign _1447 = ~ PHASE_17;
    assign write_enable_75 = _1406 & _1447;
    assign _1451 = write_enable_75 | read_enable_61;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_36
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1451), .regcea(vdd), .wea(write_enable_75), .addra(address_75), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_60), .regceb(vdd), .web(write_enable_74), .addrb(address_74), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1458[131:131]), .sbiterrb(_1458[130:130]), .doutb(_1458[129:66]), .dbiterra(_1458[65:65]), .sbiterra(_1458[64:64]), .douta(_1458[63:0]) );
    assign _1459 = _1458[63:0];
    assign _1439 = _172[11:11];
    assign _1438 = _172[10:10];
    assign _1437 = _172[9:9];
    assign _1436 = _172[8:8];
    assign _1435 = _172[7:7];
    assign _1434 = _172[6:6];
    assign _1433 = _172[5:5];
    assign _1432 = _172[4:4];
    assign _1431 = _172[3:3];
    assign _1430 = _172[2:2];
    assign _1429 = _172[1:1];
    assign _1428 = _172[0:0];
    assign _1440 = { _1428, _1429, _1430, _1431, _1432, _1433, _1434, _1435, _1436, _1437, _1438, _1439 };
    assign address_76 = PHASE_17 ? _1441 : _1440;
    assign _1425 = ~ PHASE_17;
    assign read_enable_62 = _102 & _1425;
    assign data_73 = wr_d1;
    assign _1422 = _137[11:11];
    assign _1421 = _137[10:10];
    assign _1420 = _137[9:9];
    assign _1419 = _137[8:8];
    assign _1418 = _137[7:7];
    assign _1417 = _137[6:6];
    assign _1416 = _137[5:5];
    assign _1415 = _137[4:4];
    assign _1414 = _137[3:3];
    assign _1413 = _137[2:2];
    assign _1412 = _137[1:1];
    assign _1411 = _137[0:0];
    assign _1423 = { _1411, _1412, _1413, _1414, _1415, _1416, _1417, _1418, _1419, _1420, _1421, _1422 };
    assign address_77 = PHASE_17 ? _60 : _1423;
    assign _1408 = ~ PHASE_17;
    assign read_enable_63 = _102 & _1408;
    assign _1406 = _62[1:1];
    assign write_enable_77 = _1406 & PHASE_17;
    assign _1410 = write_enable_77 | read_enable_63;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_37
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1410), .regcea(vdd), .wea(write_enable_77), .addra(address_77), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_62), .regceb(vdd), .web(write_enable_76), .addrb(address_76), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1445[131:131]), .sbiterrb(_1445[130:130]), .doutb(_1445[129:66]), .dbiterra(_1445[65:65]), .sbiterra(_1445[64:64]), .douta(_1445[63:0]) );
    assign _1446 = _1445[63:0];
    assign _1367 = ~ PHASE_17;
    assign _51 = _1367;
    always @(posedge _84) begin
        if (_82)
            PHASE_17 <= _1365;
        else
            if (_72)
                PHASE_17 <= _51;
    end
    assign _1460 = PHASE_17 ? _1459 : _1446;
    assign address_78 = _1391 ? _199 : _172;
    assign _1398 = ~ _1391;
    assign read_enable_64 = _102 & _1398;
    assign write_enable_78 = _1382 & _1391;
    assign _1400 = write_enable_78 | read_enable_64;
    assign address_79 = _1391 ? _164 : _137;
    assign _1393 = ~ _1391;
    assign read_enable_65 = _102 & _1393;
    assign _1391 = ~ PHASE_18;
    assign write_enable_79 = _1375 & _1391;
    assign _1395 = write_enable_79 | read_enable_65;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_38
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1395), .regcea(vdd), .wea(write_enable_79), .addra(address_79), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1400), .regceb(vdd), .web(write_enable_78), .addrb(address_78), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1403[131:131]), .sbiterrb(_1403[130:130]), .doutb(_1403[129:66]), .dbiterra(_1403[65:65]), .sbiterra(_1403[64:64]), .douta(_1403[63:0]) );
    assign _1404 = _1403[63:0];
    assign _1471 = _1470[127:64];
    assign data_75 = _1471;
    assign address_80 = PHASE_18 ? _199 : _172;
    assign _1384 = ~ PHASE_18;
    assign read_enable_66 = _102 & _1384;
    assign _1381 = ~ _130;
    assign _1382 = _129 & _1381;
    assign write_enable_80 = _1382 & PHASE_18;
    assign _1386 = write_enable_80 | read_enable_66;
    assign address_81 = PHASE_18 ? _164 : _137;
    assign _1377 = ~ PHASE_18;
    assign read_enable_67 = _102 & _1377;
    assign _1374 = ~ _130;
    assign _1375 = _129 & _1374;
    assign write_enable_81 = _1375 & PHASE_18;
    assign _1379 = write_enable_81 | read_enable_67;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_39
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1379), .regcea(vdd), .wea(write_enable_81), .addra(address_81), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1386), .regceb(vdd), .web(write_enable_80), .addrb(address_80), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1389[131:131]), .sbiterrb(_1389[130:130]), .doutb(_1389[129:66]), .dbiterra(_1389[65:65]), .sbiterra(_1389[64:64]), .douta(_1389[63:0]) );
    assign _1390 = _1389[63:0];
    assign _1472 = ~ PHASE_18;
    assign _53 = _1472;
    always @(posedge _84) begin
        if (_82)
            PHASE_18 <= _1372;
        else
            if (_99)
                PHASE_18 <= _53;
    end
    assign q0_5 = PHASE_18 ? _1404 : _1390;
    always @(posedge _84) begin
        if (_82)
            _1370 <= _1369;
        else
            _1370 <= _92;
    end
    assign _1461 = _1370 ? _1460 : q0_5;
    dp_0
        dp_0
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1461), .d2(_1468), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1470[191:128]), .q2(_1470[127:64]), .q1(_1470[63:0]) );
    assign _1473 = _1470[63:0];
    assign data_79 = _1473;
    assign address_82 = PHASE_19 ? _164 : _68;
    assign _1537 = ~ PHASE_19;
    assign _1536 = _70[1:1];
    assign read_enable_68 = _1536 & _1537;
    always @(posedge _84) begin
        if (_82)
            _1507 <= _1506;
        else
            _1507 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1510 <= _1509;
        else
            _1510 <= _1507;
    end
    always @(posedge _84) begin
        if (_82)
            _1513 <= _1512;
        else
            _1513 <= _1510;
    end
    always @(posedge _84) begin
        if (_82)
            _1516 <= _1515;
        else
            _1516 <= _1513;
    end
    always @(posedge _84) begin
        if (_82)
            _1519 <= _1518;
        else
            _1519 <= _1516;
    end
    always @(posedge _84) begin
        if (_82)
            _1522 <= _1521;
        else
            _1522 <= _1519;
    end
    always @(posedge _84) begin
        if (_82)
            _1525 <= _1524;
        else
            _1525 <= _1522;
    end
    always @(posedge _84) begin
        if (_82)
            _1528 <= _1527;
        else
            _1528 <= _1525;
    end
    always @(posedge _84) begin
        if (_82)
            _1531 <= _1530;
        else
            _1531 <= _1528;
    end
    assign _1532 = ~ _1531;
    always @(posedge _84) begin
        if (_82)
            _1480 <= _1479;
        else
            _1480 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1483 <= _1482;
        else
            _1483 <= _1480;
    end
    always @(posedge _84) begin
        if (_82)
            _1486 <= _1485;
        else
            _1486 <= _1483;
    end
    always @(posedge _84) begin
        if (_82)
            _1489 <= _1488;
        else
            _1489 <= _1486;
    end
    always @(posedge _84) begin
        if (_82)
            _1492 <= _1491;
        else
            _1492 <= _1489;
    end
    always @(posedge _84) begin
        if (_82)
            _1495 <= _1494;
        else
            _1495 <= _1492;
    end
    always @(posedge _84) begin
        if (_82)
            _1498 <= _1497;
        else
            _1498 <= _1495;
    end
    always @(posedge _84) begin
        if (_82)
            _1501 <= _1500;
        else
            _1501 <= _1498;
    end
    always @(posedge _84) begin
        if (_82)
            _1504 <= _1503;
        else
            _1504 <= _1501;
    end
    assign _1533 = _1504 & _1532;
    assign _1534 = _129 & _1533;
    assign write_enable_82 = _1534 & PHASE_19;
    assign _1539 = write_enable_82 | read_enable_68;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_40
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1539), .regcea(vdd), .wea(write_enable_82), .addra(address_82), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_73), .regceb(vdd), .web(write_enable_73), .addrb(address_73), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1546[131:131]), .sbiterrb(_1546[130:130]), .doutb(_1546[129:66]), .dbiterra(_1546[65:65]), .sbiterra(_1546[64:64]), .douta(_1546[63:0]) );
    assign _1547 = _1546[63:0];
    assign _1477 = ~ PHASE_19;
    assign _55 = _1477;
    always @(posedge _84) begin
        if (_82)
            PHASE_19 <= _1475;
        else
            if (_72)
                PHASE_19 <= _55;
    end
    assign _1559 = PHASE_19 ? _1558 : _1547;
    assign address_83 = _1744 ? _199 : _1739;
    assign write_enable_83 = _1737 & _1744;
    assign address_84 = _1744 ? _164 : _68;
    assign _1746 = ~ _1744;
    assign read_enable_69 = _1732 & _1746;
    assign _1744 = ~ PHASE_22;
    assign write_enable_84 = _1730 & _1744;
    assign _1748 = write_enable_84 | read_enable_69;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_41
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1748), .regcea(vdd), .wea(write_enable_84), .addra(address_84), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_83), .regceb(vdd), .web(write_enable_83), .addrb(address_83), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1753[131:131]), .sbiterrb(_1753[130:130]), .doutb(_1753[129:66]), .dbiterra(_1753[65:65]), .sbiterra(_1753[64:64]), .douta(_1753[63:0]) );
    assign _1754 = _1753[63:0];
    assign address_85 = PHASE_22 ? _199 : _1739;
    assign _1737 = _129 & _1700;
    assign write_enable_85 = _1737 & PHASE_22;
    assign _292 = _91[521:518];
    assign _291 = _91[517:517];
    assign _289 = _91[513:513];
    assign _288 = _91[512:449];
    assign _287 = _91[448:385];
    assign _286 = _91[384:321];
    assign _285 = _91[320:257];
    assign _284 = _91[256:193];
    assign _283 = _91[192:129];
    assign _282 = _91[128:65];
    assign _1662 = _1654[129:66];
    assign _1661 = _1641[129:66];
    assign _1663 = PHASE_20 ? _1662 : _1661;
    assign _1659 = _1599[129:66];
    assign _1658 = _1585[129:66];
    assign q1_6 = PHASE_21 ? _1659 : _1658;
    assign _1664 = _1566 ? _1663 : q1_6;
    assign address_86 = _1643 ? _1637 : _1636;
    assign _1649 = ~ _1643;
    assign read_enable_70 = _102 & _1649;
    assign address_87 = _1643 ? _60 : _1619;
    assign _1645 = ~ _1643;
    assign read_enable_71 = _102 & _1645;
    assign _1643 = ~ PHASE_20;
    assign write_enable_87 = _1602 & _1643;
    assign _1647 = write_enable_87 | read_enable_71;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_42
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1647), .regcea(vdd), .wea(write_enable_87), .addra(address_87), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_70), .regceb(vdd), .web(write_enable_86), .addrb(address_86), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1654[131:131]), .sbiterrb(_1654[130:130]), .doutb(_1654[129:66]), .dbiterra(_1654[65:65]), .sbiterra(_1654[64:64]), .douta(_1654[63:0]) );
    assign _1655 = _1654[63:0];
    assign _1635 = _172[11:11];
    assign _1634 = _172[10:10];
    assign _1633 = _172[9:9];
    assign _1632 = _172[8:8];
    assign _1631 = _172[7:7];
    assign _1630 = _172[6:6];
    assign _1629 = _172[5:5];
    assign _1628 = _172[4:4];
    assign _1627 = _172[3:3];
    assign _1626 = _172[2:2];
    assign _1625 = _172[1:1];
    assign _1624 = _172[0:0];
    assign _1636 = { _1624, _1625, _1626, _1627, _1628, _1629, _1630, _1631, _1632, _1633, _1634, _1635 };
    assign address_88 = PHASE_20 ? _1637 : _1636;
    assign _1621 = ~ PHASE_20;
    assign read_enable_72 = _102 & _1621;
    assign data_85 = wr_d0;
    assign _60 = wr_addr;
    assign _1618 = _137[11:11];
    assign _1617 = _137[10:10];
    assign _1616 = _137[9:9];
    assign _1615 = _137[8:8];
    assign _1614 = _137[7:7];
    assign _1613 = _137[6:6];
    assign _1612 = _137[5:5];
    assign _1611 = _137[4:4];
    assign _1610 = _137[3:3];
    assign _1609 = _137[2:2];
    assign _1608 = _137[1:1];
    assign _1607 = _137[0:0];
    assign _1619 = { _1607, _1608, _1609, _1610, _1611, _1612, _1613, _1614, _1615, _1616, _1617, _1618 };
    assign address_89 = PHASE_20 ? _60 : _1619;
    assign _1604 = ~ PHASE_20;
    assign read_enable_73 = _102 & _1604;
    assign _62 = wr_en;
    assign _1602 = _62[0:0];
    assign write_enable_89 = _1602 & PHASE_20;
    assign _1606 = write_enable_89 | read_enable_73;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_43
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1606), .regcea(vdd), .wea(write_enable_89), .addra(address_89), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_72), .regceb(vdd), .web(write_enable_88), .addrb(address_88), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1641[131:131]), .sbiterrb(_1641[130:130]), .doutb(_1641[129:66]), .dbiterra(_1641[65:65]), .sbiterra(_1641[64:64]), .douta(_1641[63:0]) );
    assign _1642 = _1641[63:0];
    assign _1563 = ~ PHASE_20;
    assign _63 = _1563;
    always @(posedge _84) begin
        if (_82)
            PHASE_20 <= _1561;
        else
            if (_72)
                PHASE_20 <= _63;
    end
    assign _1656 = PHASE_20 ? _1655 : _1642;
    assign address_90 = _1587 ? _199 : _172;
    assign _1594 = ~ _1587;
    assign read_enable_74 = _102 & _1594;
    assign write_enable_90 = _1578 & _1587;
    assign _1596 = write_enable_90 | read_enable_74;
    assign address_91 = _1587 ? _164 : _137;
    assign _1589 = ~ _1587;
    assign read_enable_75 = _102 & _1589;
    assign _1587 = ~ PHASE_21;
    assign write_enable_91 = _1571 & _1587;
    assign _1591 = write_enable_91 | read_enable_75;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_44
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1591), .regcea(vdd), .wea(write_enable_91), .addra(address_91), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1596), .regceb(vdd), .web(write_enable_90), .addrb(address_90), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1599[131:131]), .sbiterrb(_1599[130:130]), .doutb(_1599[129:66]), .dbiterra(_1599[65:65]), .sbiterra(_1599[64:64]), .douta(_1599[63:0]) );
    assign _1600 = _1599[63:0];
    assign _1667 = _1666[127:64];
    assign data_87 = _1667;
    always @(posedge _84) begin
        if (_82)
            _175 <= _174;
        else
            _175 <= _172;
    end
    always @(posedge _84) begin
        if (_82)
            _178 <= _177;
        else
            _178 <= _175;
    end
    always @(posedge _84) begin
        if (_82)
            _181 <= _180;
        else
            _181 <= _178;
    end
    always @(posedge _84) begin
        if (_82)
            _184 <= _183;
        else
            _184 <= _181;
    end
    always @(posedge _84) begin
        if (_82)
            _187 <= _186;
        else
            _187 <= _184;
    end
    always @(posedge _84) begin
        if (_82)
            _190 <= _189;
        else
            _190 <= _187;
    end
    always @(posedge _84) begin
        if (_82)
            _193 <= _192;
        else
            _193 <= _190;
    end
    always @(posedge _84) begin
        if (_82)
            _196 <= _195;
        else
            _196 <= _193;
    end
    always @(posedge _84) begin
        if (_82)
            _199 <= _198;
        else
            _199 <= _196;
    end
    assign _172 = _91[64:53];
    assign address_92 = PHASE_21 ? _199 : _172;
    assign _1580 = ~ PHASE_21;
    assign read_enable_76 = _102 & _1580;
    assign _1577 = ~ _130;
    assign _1578 = _129 & _1577;
    assign write_enable_92 = _1578 & PHASE_21;
    assign _1582 = write_enable_92 | read_enable_76;
    assign address_93 = PHASE_21 ? _164 : _137;
    assign _1573 = ~ PHASE_21;
    assign read_enable_77 = _102 & _1573;
    assign _1570 = ~ _130;
    assign _1571 = _129 & _1570;
    assign write_enable_93 = _1571 & PHASE_21;
    assign _1575 = write_enable_93 | read_enable_77;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_45
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1575), .regcea(vdd), .wea(write_enable_93), .addra(address_93), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1582), .regceb(vdd), .web(write_enable_92), .addrb(address_92), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1585[131:131]), .sbiterrb(_1585[130:130]), .doutb(_1585[129:66]), .dbiterra(_1585[65:65]), .sbiterra(_1585[64:64]), .douta(_1585[63:0]) );
    assign _1586 = _1585[63:0];
    assign _99 = _91[523:523];
    assign _1668 = ~ PHASE_21;
    assign _65 = _1668;
    always @(posedge _84) begin
        if (_82)
            PHASE_21 <= _1568;
        else
            if (_99)
                PHASE_21 <= _65;
    end
    assign q0_6 = PHASE_21 ? _1600 : _1586;
    assign _92 = _91[514:514];
    always @(posedge _84) begin
        if (_82)
            _1566 <= _1565;
        else
            _1566 <= _92;
    end
    assign _1657 = _1566 ? _1656 : q0_6;
    dp
        dp
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1657), .d2(_1664), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1666[191:128]), .q2(_1666[127:64]), .q1(_1666[63:0]) );
    assign _1669 = _1666[63:0];
    assign data_91 = _1669;
    assign _137 = _91[52:41];
    always @(posedge _84) begin
        if (_82)
            _140 <= _139;
        else
            _140 <= _137;
    end
    always @(posedge _84) begin
        if (_82)
            _143 <= _142;
        else
            _143 <= _140;
    end
    always @(posedge _84) begin
        if (_82)
            _146 <= _145;
        else
            _146 <= _143;
    end
    always @(posedge _84) begin
        if (_82)
            _149 <= _148;
        else
            _149 <= _146;
    end
    always @(posedge _84) begin
        if (_82)
            _152 <= _151;
        else
            _152 <= _149;
    end
    always @(posedge _84) begin
        if (_82)
            _155 <= _154;
        else
            _155 <= _152;
    end
    always @(posedge _84) begin
        if (_82)
            _158 <= _157;
        else
            _158 <= _155;
    end
    always @(posedge _84) begin
        if (_82)
            _161 <= _160;
        else
            _161 <= _158;
    end
    always @(posedge _84) begin
        if (_82)
            _164 <= _163;
        else
            _164 <= _161;
    end
    assign _68 = rd_addr;
    assign address_94 = PHASE_22 ? _164 : _68;
    assign _1733 = ~ PHASE_22;
    assign _70 = rd_en;
    assign _1732 = _70[0:0];
    assign read_enable_78 = _1732 & _1733;
    assign _290 = _91[516:516];
    always @(posedge _84) begin
        if (_82)
            _1703 <= _1702;
        else
            _1703 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1706 <= _1705;
        else
            _1706 <= _1703;
    end
    always @(posedge _84) begin
        if (_82)
            _1709 <= _1708;
        else
            _1709 <= _1706;
    end
    always @(posedge _84) begin
        if (_82)
            _1712 <= _1711;
        else
            _1712 <= _1709;
    end
    always @(posedge _84) begin
        if (_82)
            _1715 <= _1714;
        else
            _1715 <= _1712;
    end
    always @(posedge _84) begin
        if (_82)
            _1718 <= _1717;
        else
            _1718 <= _1715;
    end
    always @(posedge _84) begin
        if (_82)
            _1721 <= _1720;
        else
            _1721 <= _1718;
    end
    always @(posedge _84) begin
        if (_82)
            _1724 <= _1723;
        else
            _1724 <= _1721;
    end
    always @(posedge _84) begin
        if (_82)
            _1727 <= _1726;
        else
            _1727 <= _1724;
    end
    assign _1728 = ~ _1727;
    assign _130 = _91[515:515];
    always @(posedge _84) begin
        if (_82)
            _1676 <= _1675;
        else
            _1676 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1679 <= _1678;
        else
            _1679 <= _1676;
    end
    always @(posedge _84) begin
        if (_82)
            _1682 <= _1681;
        else
            _1682 <= _1679;
    end
    always @(posedge _84) begin
        if (_82)
            _1685 <= _1684;
        else
            _1685 <= _1682;
    end
    always @(posedge _84) begin
        if (_82)
            _1688 <= _1687;
        else
            _1688 <= _1685;
    end
    always @(posedge _84) begin
        if (_82)
            _1691 <= _1690;
        else
            _1691 <= _1688;
    end
    always @(posedge _84) begin
        if (_82)
            _1694 <= _1693;
        else
            _1694 <= _1691;
    end
    always @(posedge _84) begin
        if (_82)
            _1697 <= _1696;
        else
            _1697 <= _1694;
    end
    always @(posedge _84) begin
        if (_82)
            _1700 <= _1699;
        else
            _1700 <= _1697;
    end
    assign _1729 = _1700 & _1728;
    assign _102 = _91[522:522];
    always @(posedge _84) begin
        if (_82)
            _105 <= _104;
        else
            _105 <= _102;
    end
    always @(posedge _84) begin
        if (_82)
            _108 <= _107;
        else
            _108 <= _105;
    end
    always @(posedge _84) begin
        if (_82)
            _111 <= _110;
        else
            _111 <= _108;
    end
    always @(posedge _84) begin
        if (_82)
            _114 <= _113;
        else
            _114 <= _111;
    end
    always @(posedge _84) begin
        if (_82)
            _117 <= _116;
        else
            _117 <= _114;
    end
    always @(posedge _84) begin
        if (_82)
            _120 <= _119;
        else
            _120 <= _117;
    end
    always @(posedge _84) begin
        if (_82)
            _123 <= _122;
        else
            _123 <= _120;
    end
    always @(posedge _84) begin
        if (_82)
            _126 <= _125;
        else
            _126 <= _123;
    end
    always @(posedge _84) begin
        if (_82)
            _129 <= _128;
        else
            _129 <= _126;
    end
    assign _1730 = _129 & _1729;
    assign write_enable_94 = _1730 & PHASE_22;
    assign _1735 = write_enable_94 | read_enable_78;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_46
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1735), .regcea(vdd), .wea(write_enable_94), .addra(address_94), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_85), .regceb(vdd), .web(write_enable_85), .addrb(address_85), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1742[131:131]), .sbiterrb(_1742[130:130]), .doutb(_1742[129:66]), .dbiterra(_1742[65:65]), .sbiterra(_1742[64:64]), .douta(_1742[63:0]) );
    assign _1743 = _1742[63:0];
    assign _72 = flip;
    assign _1673 = ~ PHASE_22;
    assign _73 = _1673;
    always @(posedge _84) begin
        if (_82)
            PHASE_22 <= _1671;
        else
            if (_72)
                PHASE_22 <= _73;
    end
    assign _1755 = PHASE_22 ? _1754 : _1743;
    assign _76 = first_4step_pass;
    assign _78 = first_iter;
    assign _80 = start;
    assign _82 = clear;
    assign _84 = clock;
    ctrl
        ctrl
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .first_4step_pass(_76), .flip(_91[523:523]), .read_write_enable(_91[522:522]), .index(_91[521:518]), .valid(_91[517:517]), .twiddle_stage(_91[516:516]), .last_stage(_91[515:515]), .first_stage(_91[514:514]), .start_twiddles(_91[513:513]), .omegas6(_91[512:449]), .omegas5(_91[448:385]), .omegas4(_91[384:321]), .omegas3(_91[320:257]), .omegas2(_91[256:193]), .omegas1(_91[192:129]), .omegas0(_91[128:65]), .addr2(_91[64:53]), .addr1(_91[52:41]), .m(_91[40:29]), .k(_91[28:17]), .j(_91[16:5]), .i(_91[4:1]), .done_(_91[0:0]) );
    assign _1756 = _91[0:0];

    /* aliases */
    assign data_0 = data;
    assign data_2 = data_1;
    assign data_4 = data_3;
    assign data_5 = data_3;
    assign data_6 = data_3;
    assign data_8 = data_7;
    assign data_9 = data_7;
    assign data_10 = data_7;
    assign data_12 = data_11;
    assign data_14 = data_13;
    assign data_16 = data_15;
    assign data_17 = data_15;
    assign data_18 = data_15;
    assign data_20 = data_19;
    assign data_21 = data_19;
    assign data_22 = data_19;
    assign data_24 = data_23;
    assign data_26 = data_25;
    assign data_28 = data_27;
    assign data_29 = data_27;
    assign data_30 = data_27;
    assign data_32 = data_31;
    assign data_33 = data_31;
    assign data_34 = data_31;
    assign data_36 = data_35;
    assign data_38 = data_37;
    assign data_40 = data_39;
    assign data_41 = data_39;
    assign data_42 = data_39;
    assign data_44 = data_43;
    assign data_45 = data_43;
    assign data_46 = data_43;
    assign data_48 = data_47;
    assign data_50 = data_49;
    assign data_52 = data_51;
    assign data_53 = data_51;
    assign data_54 = data_51;
    assign data_56 = data_55;
    assign data_57 = data_55;
    assign data_58 = data_55;
    assign data_60 = data_59;
    assign data_62 = data_61;
    assign data_64 = data_63;
    assign data_65 = data_63;
    assign data_66 = data_63;
    assign data_68 = data_67;
    assign data_69 = data_67;
    assign data_70 = data_67;
    assign data_72 = data_71;
    assign data_74 = data_73;
    assign data_76 = data_75;
    assign data_77 = data_75;
    assign data_78 = data_75;
    assign data_80 = data_79;
    assign data_81 = data_79;
    assign data_82 = data_79;
    assign data_84 = data_83;
    assign data_86 = data_85;
    assign data_88 = data_87;
    assign data_89 = data_87;
    assign data_90 = data_87;
    assign data_92 = data_91;
    assign data_93 = data_91;
    assign data_94 = data_91;

    /* output assignments */
    assign done_ = _1756;
    assign rd_q0 = _1755;
    assign rd_q1 = _1559;
    assign rd_q2 = _1363;
    assign rd_q3 = _1167;
    assign rd_q4 = _971;
    assign rd_q5 = _775;
    assign rd_q6 = _579;
    assign rd_q7 = _383;

endmodule
module dp_7 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0100000001000101111010011110100001010111011001101011110100011101;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0000101011001010001100100100101101011011001100100000011011011100;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1100111100000101001110011010010101001111101000110101101001010101;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1111101111010100000111000110101110001100101010100011001100000010;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0010101111111100010110000001100000101010110111101101100011110100;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0011000010111010001011101100110101011110100100111110011101101101;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1111010100000010101011101111010100110010001100100010011001010100;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_8 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0000010100100101000010101011110010110110000000011111001101101000;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0000000010100111001011000000010010100111011101011111110001111000;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0101010110001110111110001100010010001010101000010011001111000110;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0110110010110000111011001100000000010111101011101101100010111100;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0111110100110000011011110001001011110110100001101100011000110001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1111011001111000001001110011001110101011000101110000100110010000;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1000000110000100011111010011111110001100111000110111011110101010;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_9 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1100001011100100110011000100001001100010000010000101000110100011;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0101100000001101011100101110110101101100101000101100101011001111;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0001100100000101011100000100110001000100110010001101110010111010;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1100111100000101001110011010010101001111101000110101101001010101;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1101100000000001010001101110001110101111011110010110111001001011;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1100101111011100100111001010001111010111100111010001110111111011;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1100110100011111000010100001011101001011100011010101101111000110;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_10 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1011010110101101000000101101111100111100001110110110000100100100;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0110100101101111110010001001101110011101101001011110000011100001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0000110011111011010001010110001011100101111101011000011111100101;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1101101000101011101011101011110001010010100001010000110110101000;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1100001001011111000111001110000000001100100011011001101101100111;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1100100111010010110100011100111101011011010100100100011110000101;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1111010111110011111101100110101110011110000000010111000110010101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_11 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0110001110111000011110101101110010111010001011110110000001100110;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0000000110011111011011110111001101111001110110010011010011110001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0101100000001101011100101110110101101100101000101100101011001111;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0000101011001010001100100100101101011011001100100000011011011100;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0110110010110000111011001100000000010111101011101101100010111100;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0010101111111100010110000001100000101010110111101101100011110100;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1110100111111101110111001000100000111011101101000001000000101001;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_12 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0100000001110001000111111100111100100111011110111011010011010110;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0010111110010100110000110000001100100101110011011100011011100111;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0011101100101111111010001010011101110000101100100110000011010001;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1000011011100101001000010011100100111101111001011101100010110100;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0001001110110001100110001111101111010100011111111100000011111001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0011101010000111001111101001111000100100000111000010101101000010;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0011011000110010000010101111100100011101101001111100011001110011;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_13 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1000000110101110110111001110001000000110110000010101010010110101;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0110001110111000011110101101110010111010001011110110000001100110;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1100001011100100110011000100001001100010000010000101000110100011;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0100000001000101111010011110100001010111011001101011110100011101;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0010101001001000011111010001011101101011111100000111111100100010;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0000110110101000001001111111111011110100101101110111101011101101;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0000101000011000111111101100011111011101011101011111000010111001;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_14 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0101110100110000000100110101011101000010111111000111010000001011;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0100000110110111010100110011011100010101000101100000000101100101;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1011001001111110010011100100101001101101101011111111101111011111;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0101100000001101011100101110110101101100101000101100101011001111;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0101010110001110111110001100010010001010101000010011001111000110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1101100000000001010001101110001110101111011110010110111001001011;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0010000100100010111110011011000001011110111001100011000101100111;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module parallel_cores_0 (
    wr_d7,
    wr_d6,
    wr_d5,
    wr_d4,
    wr_d3,
    wr_d2,
    wr_d1,
    wr_d0,
    wr_addr,
    wr_en,
    rd_addr,
    rd_en,
    flip,
    first_4step_pass,
    first_iter,
    start,
    clear,
    clock,
    done_,
    rd_q0,
    rd_q1,
    rd_q2,
    rd_q3,
    rd_q4,
    rd_q5,
    rd_q6,
    rd_q7
);

    input [63:0] wr_d7;
    input [63:0] wr_d6;
    input [63:0] wr_d5;
    input [63:0] wr_d4;
    input [63:0] wr_d3;
    input [63:0] wr_d2;
    input [63:0] wr_d1;
    input [63:0] wr_d0;
    input [11:0] wr_addr;
    input [7:0] wr_en;
    input [11:0] rd_addr;
    input [7:0] rd_en;
    input flip;
    input first_4step_pass;
    input first_iter;
    input start;
    input clear;
    input clock;
    output done_;
    output [63:0] rd_q0;
    output [63:0] rd_q1;
    output [63:0] rd_q2;
    output [63:0] rd_q3;
    output [63:0] rd_q4;
    output [63:0] rd_q5;
    output [63:0] rd_q6;
    output [63:0] rd_q7;

    /* signal declarations */
    wire [11:0] address;
    wire write_enable;
    wire [11:0] address_0;
    wire _374;
    wire read_enable;
    wire _372;
    wire write_enable_0;
    wire _376;
    wire [131:0] _381;
    wire [63:0] _382;
    wire [11:0] _367 = 12'b000000000000;
    wire [11:0] address_1;
    wire _365;
    wire write_enable_1;
    wire [63:0] _279;
    wire [63:0] _278;
    wire [63:0] _280;
    wire [63:0] _276;
    wire [63:0] _275;
    wire [63:0] q1;
    wire [63:0] _281;
    wire [11:0] address_2;
    wire write_enable_2 = 1'b0;
    wire _266;
    wire read_enable_0;
    wire [11:0] address_3;
    wire _262;
    wire read_enable_1;
    wire _260;
    wire write_enable_3;
    wire _264;
    wire [131:0] _271;
    wire [63:0] _272;
    wire [63:0] data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_0;
    wire [11:0] _254 = 12'b000000000000;
    wire _252;
    wire _251;
    wire _250;
    wire _249;
    wire _248;
    wire _247;
    wire _246;
    wire _245;
    wire _244;
    wire _243;
    wire _242;
    wire _241;
    wire [11:0] _253;
    wire [11:0] address_4;
    wire write_enable_4 = 1'b0;
    wire _238;
    wire read_enable_2;
    wire [63:0] data_1;
    wire [63:0] data_2;
    wire _235;
    wire _234;
    wire _233;
    wire _232;
    wire _231;
    wire _230;
    wire _229;
    wire _228;
    wire _227;
    wire _226;
    wire _225;
    wire _224;
    wire [11:0] _236;
    wire [11:0] address_5;
    wire _221;
    wire read_enable_3;
    wire _219;
    wire write_enable_5;
    wire _223;
    wire [131:0] _258;
    wire [63:0] _259;
    wire _87 = 1'b0;
    wire _86 = 1'b0;
    wire _89;
    wire _3;
    reg PHASE;
    wire [63:0] _273;
    wire [11:0] address_6;
    wire _211;
    wire read_enable_4;
    wire write_enable_6;
    wire _213;
    wire [11:0] address_7;
    wire _206;
    wire read_enable_5;
    wire _204;
    wire write_enable_7;
    wire _208;
    wire [131:0] _216;
    wire [63:0] _217;
    wire [63:0] _295;
    wire [63:0] data_3;
    wire [63:0] data_4;
    wire [63:0] data_5;
    wire [63:0] data_6;
    wire [11:0] address_8;
    wire _169;
    wire read_enable_6;
    wire _166;
    wire _167;
    wire write_enable_8;
    wire _171;
    wire [11:0] address_9;
    wire _134;
    wire read_enable_7;
    wire _131;
    wire _132;
    wire write_enable_9;
    wire _136;
    wire [131:0] _202;
    wire [63:0] _203;
    wire _98 = 1'b0;
    wire _97 = 1'b0;
    wire _296;
    wire _5;
    reg PHASE_0;
    wire [63:0] q0;
    wire _94 = 1'b0;
    wire _93 = 1'b0;
    reg _96;
    wire [63:0] _274;
    wire [191:0] _294;
    wire [63:0] _297;
    wire [63:0] data_7;
    wire [63:0] data_8;
    wire [63:0] data_9;
    wire [63:0] data_10;
    wire [11:0] address_10;
    wire _361;
    wire _360;
    wire read_enable_8;
    wire _354 = 1'b0;
    wire _353 = 1'b0;
    wire _351 = 1'b0;
    wire _350 = 1'b0;
    wire _348 = 1'b0;
    wire _347 = 1'b0;
    wire _345 = 1'b0;
    wire _344 = 1'b0;
    wire _342 = 1'b0;
    wire _341 = 1'b0;
    wire _339 = 1'b0;
    wire _338 = 1'b0;
    wire _336 = 1'b0;
    wire _335 = 1'b0;
    wire _333 = 1'b0;
    wire _332 = 1'b0;
    wire _330 = 1'b0;
    wire _329 = 1'b0;
    reg _331;
    reg _334;
    reg _337;
    reg _340;
    reg _343;
    reg _346;
    reg _349;
    reg _352;
    reg _355;
    wire _356;
    wire _327 = 1'b0;
    wire _326 = 1'b0;
    wire _324 = 1'b0;
    wire _323 = 1'b0;
    wire _321 = 1'b0;
    wire _320 = 1'b0;
    wire _318 = 1'b0;
    wire _317 = 1'b0;
    wire _315 = 1'b0;
    wire _314 = 1'b0;
    wire _312 = 1'b0;
    wire _311 = 1'b0;
    wire _309 = 1'b0;
    wire _308 = 1'b0;
    wire _306 = 1'b0;
    wire _305 = 1'b0;
    wire _303 = 1'b0;
    wire _302 = 1'b0;
    reg _304;
    reg _307;
    reg _310;
    reg _313;
    reg _316;
    reg _319;
    reg _322;
    reg _325;
    reg _328;
    wire _357;
    wire _358;
    wire write_enable_10;
    wire _363;
    wire [131:0] _370;
    wire [63:0] _371;
    wire _299 = 1'b0;
    wire _298 = 1'b0;
    wire _301;
    wire _7;
    reg PHASE_1;
    wire [63:0] _383;
    wire [11:0] address_11;
    wire write_enable_11;
    wire [11:0] address_12;
    wire _570;
    wire read_enable_9;
    wire _568;
    wire write_enable_12;
    wire _572;
    wire [131:0] _577;
    wire [63:0] _578;
    wire [11:0] _563 = 12'b000000000000;
    wire [11:0] address_13;
    wire _561;
    wire write_enable_13;
    wire [63:0] _486;
    wire [63:0] _485;
    wire [63:0] _487;
    wire [63:0] _483;
    wire [63:0] _482;
    wire [63:0] q1_0;
    wire [63:0] _488;
    wire [11:0] address_14;
    wire write_enable_14 = 1'b0;
    wire _473;
    wire read_enable_10;
    wire [11:0] address_15;
    wire _469;
    wire read_enable_11;
    wire _467;
    wire write_enable_15;
    wire _471;
    wire [131:0] _478;
    wire [63:0] _479;
    wire [63:0] data_11 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_12;
    wire [11:0] _461 = 12'b000000000000;
    wire _459;
    wire _458;
    wire _457;
    wire _456;
    wire _455;
    wire _454;
    wire _453;
    wire _452;
    wire _451;
    wire _450;
    wire _449;
    wire _448;
    wire [11:0] _460;
    wire [11:0] address_16;
    wire write_enable_16 = 1'b0;
    wire _445;
    wire read_enable_12;
    wire [63:0] data_13;
    wire [63:0] data_14;
    wire _442;
    wire _441;
    wire _440;
    wire _439;
    wire _438;
    wire _437;
    wire _436;
    wire _435;
    wire _434;
    wire _433;
    wire _432;
    wire _431;
    wire [11:0] _443;
    wire [11:0] address_17;
    wire _428;
    wire read_enable_13;
    wire _426;
    wire write_enable_17;
    wire _430;
    wire [131:0] _465;
    wire [63:0] _466;
    wire _385 = 1'b0;
    wire _384 = 1'b0;
    wire _387;
    wire _11;
    reg PHASE_2;
    wire [63:0] _480;
    wire [11:0] address_18;
    wire _418;
    wire read_enable_14;
    wire write_enable_18;
    wire _420;
    wire [11:0] address_19;
    wire _413;
    wire read_enable_15;
    wire _411;
    wire write_enable_19;
    wire _415;
    wire [131:0] _423;
    wire [63:0] _424;
    wire [63:0] _491;
    wire [63:0] data_15;
    wire [63:0] data_16;
    wire [63:0] data_17;
    wire [63:0] data_18;
    wire [11:0] address_20;
    wire _404;
    wire read_enable_16;
    wire _401;
    wire _402;
    wire write_enable_20;
    wire _406;
    wire [11:0] address_21;
    wire _397;
    wire read_enable_17;
    wire _394;
    wire _395;
    wire write_enable_21;
    wire _399;
    wire [131:0] _409;
    wire [63:0] _410;
    wire _392 = 1'b0;
    wire _391 = 1'b0;
    wire _492;
    wire _13;
    reg PHASE_3;
    wire [63:0] q0_0;
    wire _389 = 1'b0;
    wire _388 = 1'b0;
    reg _390;
    wire [63:0] _481;
    wire [191:0] _490;
    wire [63:0] _493;
    wire [63:0] data_19;
    wire [63:0] data_20;
    wire [63:0] data_21;
    wire [63:0] data_22;
    wire [11:0] address_22;
    wire _557;
    wire _556;
    wire read_enable_18;
    wire _550 = 1'b0;
    wire _549 = 1'b0;
    wire _547 = 1'b0;
    wire _546 = 1'b0;
    wire _544 = 1'b0;
    wire _543 = 1'b0;
    wire _541 = 1'b0;
    wire _540 = 1'b0;
    wire _538 = 1'b0;
    wire _537 = 1'b0;
    wire _535 = 1'b0;
    wire _534 = 1'b0;
    wire _532 = 1'b0;
    wire _531 = 1'b0;
    wire _529 = 1'b0;
    wire _528 = 1'b0;
    wire _526 = 1'b0;
    wire _525 = 1'b0;
    reg _527;
    reg _530;
    reg _533;
    reg _536;
    reg _539;
    reg _542;
    reg _545;
    reg _548;
    reg _551;
    wire _552;
    wire _523 = 1'b0;
    wire _522 = 1'b0;
    wire _520 = 1'b0;
    wire _519 = 1'b0;
    wire _517 = 1'b0;
    wire _516 = 1'b0;
    wire _514 = 1'b0;
    wire _513 = 1'b0;
    wire _511 = 1'b0;
    wire _510 = 1'b0;
    wire _508 = 1'b0;
    wire _507 = 1'b0;
    wire _505 = 1'b0;
    wire _504 = 1'b0;
    wire _502 = 1'b0;
    wire _501 = 1'b0;
    wire _499 = 1'b0;
    wire _498 = 1'b0;
    reg _500;
    reg _503;
    reg _506;
    reg _509;
    reg _512;
    reg _515;
    reg _518;
    reg _521;
    reg _524;
    wire _553;
    wire _554;
    wire write_enable_22;
    wire _559;
    wire [131:0] _566;
    wire [63:0] _567;
    wire _495 = 1'b0;
    wire _494 = 1'b0;
    wire _497;
    wire _15;
    reg PHASE_4;
    wire [63:0] _579;
    wire [11:0] address_23;
    wire write_enable_23;
    wire [11:0] address_24;
    wire _766;
    wire read_enable_19;
    wire _764;
    wire write_enable_24;
    wire _768;
    wire [131:0] _773;
    wire [63:0] _774;
    wire [11:0] _759 = 12'b000000000000;
    wire [11:0] address_25;
    wire _757;
    wire write_enable_25;
    wire [63:0] _682;
    wire [63:0] _681;
    wire [63:0] _683;
    wire [63:0] _679;
    wire [63:0] _678;
    wire [63:0] q1_1;
    wire [63:0] _684;
    wire [11:0] address_26;
    wire write_enable_26 = 1'b0;
    wire _669;
    wire read_enable_20;
    wire [11:0] address_27;
    wire _665;
    wire read_enable_21;
    wire _663;
    wire write_enable_27;
    wire _667;
    wire [131:0] _674;
    wire [63:0] _675;
    wire [63:0] data_23 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_24;
    wire [11:0] _657 = 12'b000000000000;
    wire _655;
    wire _654;
    wire _653;
    wire _652;
    wire _651;
    wire _650;
    wire _649;
    wire _648;
    wire _647;
    wire _646;
    wire _645;
    wire _644;
    wire [11:0] _656;
    wire [11:0] address_28;
    wire write_enable_28 = 1'b0;
    wire _641;
    wire read_enable_22;
    wire [63:0] data_25;
    wire [63:0] data_26;
    wire _638;
    wire _637;
    wire _636;
    wire _635;
    wire _634;
    wire _633;
    wire _632;
    wire _631;
    wire _630;
    wire _629;
    wire _628;
    wire _627;
    wire [11:0] _639;
    wire [11:0] address_29;
    wire _624;
    wire read_enable_23;
    wire _622;
    wire write_enable_29;
    wire _626;
    wire [131:0] _661;
    wire [63:0] _662;
    wire _581 = 1'b0;
    wire _580 = 1'b0;
    wire _583;
    wire _19;
    reg PHASE_5;
    wire [63:0] _676;
    wire [11:0] address_30;
    wire _614;
    wire read_enable_24;
    wire write_enable_30;
    wire _616;
    wire [11:0] address_31;
    wire _609;
    wire read_enable_25;
    wire _607;
    wire write_enable_31;
    wire _611;
    wire [131:0] _619;
    wire [63:0] _620;
    wire [63:0] _687;
    wire [63:0] data_27;
    wire [63:0] data_28;
    wire [63:0] data_29;
    wire [63:0] data_30;
    wire [11:0] address_32;
    wire _600;
    wire read_enable_26;
    wire _597;
    wire _598;
    wire write_enable_32;
    wire _602;
    wire [11:0] address_33;
    wire _593;
    wire read_enable_27;
    wire _590;
    wire _591;
    wire write_enable_33;
    wire _595;
    wire [131:0] _605;
    wire [63:0] _606;
    wire _588 = 1'b0;
    wire _587 = 1'b0;
    wire _688;
    wire _21;
    reg PHASE_6;
    wire [63:0] q0_1;
    wire _585 = 1'b0;
    wire _584 = 1'b0;
    reg _586;
    wire [63:0] _677;
    wire [191:0] _686;
    wire [63:0] _689;
    wire [63:0] data_31;
    wire [63:0] data_32;
    wire [63:0] data_33;
    wire [63:0] data_34;
    wire [11:0] address_34;
    wire _753;
    wire _752;
    wire read_enable_28;
    wire _746 = 1'b0;
    wire _745 = 1'b0;
    wire _743 = 1'b0;
    wire _742 = 1'b0;
    wire _740 = 1'b0;
    wire _739 = 1'b0;
    wire _737 = 1'b0;
    wire _736 = 1'b0;
    wire _734 = 1'b0;
    wire _733 = 1'b0;
    wire _731 = 1'b0;
    wire _730 = 1'b0;
    wire _728 = 1'b0;
    wire _727 = 1'b0;
    wire _725 = 1'b0;
    wire _724 = 1'b0;
    wire _722 = 1'b0;
    wire _721 = 1'b0;
    reg _723;
    reg _726;
    reg _729;
    reg _732;
    reg _735;
    reg _738;
    reg _741;
    reg _744;
    reg _747;
    wire _748;
    wire _719 = 1'b0;
    wire _718 = 1'b0;
    wire _716 = 1'b0;
    wire _715 = 1'b0;
    wire _713 = 1'b0;
    wire _712 = 1'b0;
    wire _710 = 1'b0;
    wire _709 = 1'b0;
    wire _707 = 1'b0;
    wire _706 = 1'b0;
    wire _704 = 1'b0;
    wire _703 = 1'b0;
    wire _701 = 1'b0;
    wire _700 = 1'b0;
    wire _698 = 1'b0;
    wire _697 = 1'b0;
    wire _695 = 1'b0;
    wire _694 = 1'b0;
    reg _696;
    reg _699;
    reg _702;
    reg _705;
    reg _708;
    reg _711;
    reg _714;
    reg _717;
    reg _720;
    wire _749;
    wire _750;
    wire write_enable_34;
    wire _755;
    wire [131:0] _762;
    wire [63:0] _763;
    wire _691 = 1'b0;
    wire _690 = 1'b0;
    wire _693;
    wire _23;
    reg PHASE_7;
    wire [63:0] _775;
    wire [11:0] address_35;
    wire write_enable_35;
    wire [11:0] address_36;
    wire _962;
    wire read_enable_29;
    wire _960;
    wire write_enable_36;
    wire _964;
    wire [131:0] _969;
    wire [63:0] _970;
    wire [11:0] _955 = 12'b000000000000;
    wire [11:0] address_37;
    wire _953;
    wire write_enable_37;
    wire [63:0] _878;
    wire [63:0] _877;
    wire [63:0] _879;
    wire [63:0] _875;
    wire [63:0] _874;
    wire [63:0] q1_2;
    wire [63:0] _880;
    wire [11:0] address_38;
    wire write_enable_38 = 1'b0;
    wire _865;
    wire read_enable_30;
    wire [11:0] address_39;
    wire _861;
    wire read_enable_31;
    wire _859;
    wire write_enable_39;
    wire _863;
    wire [131:0] _870;
    wire [63:0] _871;
    wire [63:0] data_35 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_36;
    wire [11:0] _853 = 12'b000000000000;
    wire _851;
    wire _850;
    wire _849;
    wire _848;
    wire _847;
    wire _846;
    wire _845;
    wire _844;
    wire _843;
    wire _842;
    wire _841;
    wire _840;
    wire [11:0] _852;
    wire [11:0] address_40;
    wire write_enable_40 = 1'b0;
    wire _837;
    wire read_enable_32;
    wire [63:0] data_37;
    wire [63:0] data_38;
    wire _834;
    wire _833;
    wire _832;
    wire _831;
    wire _830;
    wire _829;
    wire _828;
    wire _827;
    wire _826;
    wire _825;
    wire _824;
    wire _823;
    wire [11:0] _835;
    wire [11:0] address_41;
    wire _820;
    wire read_enable_33;
    wire _818;
    wire write_enable_41;
    wire _822;
    wire [131:0] _857;
    wire [63:0] _858;
    wire _777 = 1'b0;
    wire _776 = 1'b0;
    wire _779;
    wire _27;
    reg PHASE_8;
    wire [63:0] _872;
    wire [11:0] address_42;
    wire _810;
    wire read_enable_34;
    wire write_enable_42;
    wire _812;
    wire [11:0] address_43;
    wire _805;
    wire read_enable_35;
    wire _803;
    wire write_enable_43;
    wire _807;
    wire [131:0] _815;
    wire [63:0] _816;
    wire [63:0] _883;
    wire [63:0] data_39;
    wire [63:0] data_40;
    wire [63:0] data_41;
    wire [63:0] data_42;
    wire [11:0] address_44;
    wire _796;
    wire read_enable_36;
    wire _793;
    wire _794;
    wire write_enable_44;
    wire _798;
    wire [11:0] address_45;
    wire _789;
    wire read_enable_37;
    wire _786;
    wire _787;
    wire write_enable_45;
    wire _791;
    wire [131:0] _801;
    wire [63:0] _802;
    wire _784 = 1'b0;
    wire _783 = 1'b0;
    wire _884;
    wire _29;
    reg PHASE_9;
    wire [63:0] q0_2;
    wire _781 = 1'b0;
    wire _780 = 1'b0;
    reg _782;
    wire [63:0] _873;
    wire [191:0] _882;
    wire [63:0] _885;
    wire [63:0] data_43;
    wire [63:0] data_44;
    wire [63:0] data_45;
    wire [63:0] data_46;
    wire [11:0] address_46;
    wire _949;
    wire _948;
    wire read_enable_38;
    wire _942 = 1'b0;
    wire _941 = 1'b0;
    wire _939 = 1'b0;
    wire _938 = 1'b0;
    wire _936 = 1'b0;
    wire _935 = 1'b0;
    wire _933 = 1'b0;
    wire _932 = 1'b0;
    wire _930 = 1'b0;
    wire _929 = 1'b0;
    wire _927 = 1'b0;
    wire _926 = 1'b0;
    wire _924 = 1'b0;
    wire _923 = 1'b0;
    wire _921 = 1'b0;
    wire _920 = 1'b0;
    wire _918 = 1'b0;
    wire _917 = 1'b0;
    reg _919;
    reg _922;
    reg _925;
    reg _928;
    reg _931;
    reg _934;
    reg _937;
    reg _940;
    reg _943;
    wire _944;
    wire _915 = 1'b0;
    wire _914 = 1'b0;
    wire _912 = 1'b0;
    wire _911 = 1'b0;
    wire _909 = 1'b0;
    wire _908 = 1'b0;
    wire _906 = 1'b0;
    wire _905 = 1'b0;
    wire _903 = 1'b0;
    wire _902 = 1'b0;
    wire _900 = 1'b0;
    wire _899 = 1'b0;
    wire _897 = 1'b0;
    wire _896 = 1'b0;
    wire _894 = 1'b0;
    wire _893 = 1'b0;
    wire _891 = 1'b0;
    wire _890 = 1'b0;
    reg _892;
    reg _895;
    reg _898;
    reg _901;
    reg _904;
    reg _907;
    reg _910;
    reg _913;
    reg _916;
    wire _945;
    wire _946;
    wire write_enable_46;
    wire _951;
    wire [131:0] _958;
    wire [63:0] _959;
    wire _887 = 1'b0;
    wire _886 = 1'b0;
    wire _889;
    wire _31;
    reg PHASE_10;
    wire [63:0] _971;
    wire [11:0] address_47;
    wire write_enable_47;
    wire [11:0] address_48;
    wire _1158;
    wire read_enable_39;
    wire _1156;
    wire write_enable_48;
    wire _1160;
    wire [131:0] _1165;
    wire [63:0] _1166;
    wire [11:0] _1151 = 12'b000000000000;
    wire [11:0] address_49;
    wire _1149;
    wire write_enable_49;
    wire [63:0] _1074;
    wire [63:0] _1073;
    wire [63:0] _1075;
    wire [63:0] _1071;
    wire [63:0] _1070;
    wire [63:0] q1_3;
    wire [63:0] _1076;
    wire [11:0] address_50;
    wire write_enable_50 = 1'b0;
    wire _1061;
    wire read_enable_40;
    wire [11:0] address_51;
    wire _1057;
    wire read_enable_41;
    wire _1055;
    wire write_enable_51;
    wire _1059;
    wire [131:0] _1066;
    wire [63:0] _1067;
    wire [63:0] data_47 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_48;
    wire [11:0] _1049 = 12'b000000000000;
    wire _1047;
    wire _1046;
    wire _1045;
    wire _1044;
    wire _1043;
    wire _1042;
    wire _1041;
    wire _1040;
    wire _1039;
    wire _1038;
    wire _1037;
    wire _1036;
    wire [11:0] _1048;
    wire [11:0] address_52;
    wire write_enable_52 = 1'b0;
    wire _1033;
    wire read_enable_42;
    wire [63:0] data_49;
    wire [63:0] data_50;
    wire _1030;
    wire _1029;
    wire _1028;
    wire _1027;
    wire _1026;
    wire _1025;
    wire _1024;
    wire _1023;
    wire _1022;
    wire _1021;
    wire _1020;
    wire _1019;
    wire [11:0] _1031;
    wire [11:0] address_53;
    wire _1016;
    wire read_enable_43;
    wire _1014;
    wire write_enable_53;
    wire _1018;
    wire [131:0] _1053;
    wire [63:0] _1054;
    wire _973 = 1'b0;
    wire _972 = 1'b0;
    wire _975;
    wire _35;
    reg PHASE_11;
    wire [63:0] _1068;
    wire [11:0] address_54;
    wire _1006;
    wire read_enable_44;
    wire write_enable_54;
    wire _1008;
    wire [11:0] address_55;
    wire _1001;
    wire read_enable_45;
    wire _999;
    wire write_enable_55;
    wire _1003;
    wire [131:0] _1011;
    wire [63:0] _1012;
    wire [63:0] _1079;
    wire [63:0] data_51;
    wire [63:0] data_52;
    wire [63:0] data_53;
    wire [63:0] data_54;
    wire [11:0] address_56;
    wire _992;
    wire read_enable_46;
    wire _989;
    wire _990;
    wire write_enable_56;
    wire _994;
    wire [11:0] address_57;
    wire _985;
    wire read_enable_47;
    wire _982;
    wire _983;
    wire write_enable_57;
    wire _987;
    wire [131:0] _997;
    wire [63:0] _998;
    wire _980 = 1'b0;
    wire _979 = 1'b0;
    wire _1080;
    wire _37;
    reg PHASE_12;
    wire [63:0] q0_3;
    wire _977 = 1'b0;
    wire _976 = 1'b0;
    reg _978;
    wire [63:0] _1069;
    wire [191:0] _1078;
    wire [63:0] _1081;
    wire [63:0] data_55;
    wire [63:0] data_56;
    wire [63:0] data_57;
    wire [63:0] data_58;
    wire [11:0] address_58;
    wire _1145;
    wire _1144;
    wire read_enable_48;
    wire _1138 = 1'b0;
    wire _1137 = 1'b0;
    wire _1135 = 1'b0;
    wire _1134 = 1'b0;
    wire _1132 = 1'b0;
    wire _1131 = 1'b0;
    wire _1129 = 1'b0;
    wire _1128 = 1'b0;
    wire _1126 = 1'b0;
    wire _1125 = 1'b0;
    wire _1123 = 1'b0;
    wire _1122 = 1'b0;
    wire _1120 = 1'b0;
    wire _1119 = 1'b0;
    wire _1117 = 1'b0;
    wire _1116 = 1'b0;
    wire _1114 = 1'b0;
    wire _1113 = 1'b0;
    reg _1115;
    reg _1118;
    reg _1121;
    reg _1124;
    reg _1127;
    reg _1130;
    reg _1133;
    reg _1136;
    reg _1139;
    wire _1140;
    wire _1111 = 1'b0;
    wire _1110 = 1'b0;
    wire _1108 = 1'b0;
    wire _1107 = 1'b0;
    wire _1105 = 1'b0;
    wire _1104 = 1'b0;
    wire _1102 = 1'b0;
    wire _1101 = 1'b0;
    wire _1099 = 1'b0;
    wire _1098 = 1'b0;
    wire _1096 = 1'b0;
    wire _1095 = 1'b0;
    wire _1093 = 1'b0;
    wire _1092 = 1'b0;
    wire _1090 = 1'b0;
    wire _1089 = 1'b0;
    wire _1087 = 1'b0;
    wire _1086 = 1'b0;
    reg _1088;
    reg _1091;
    reg _1094;
    reg _1097;
    reg _1100;
    reg _1103;
    reg _1106;
    reg _1109;
    reg _1112;
    wire _1141;
    wire _1142;
    wire write_enable_58;
    wire _1147;
    wire [131:0] _1154;
    wire [63:0] _1155;
    wire _1083 = 1'b0;
    wire _1082 = 1'b0;
    wire _1085;
    wire _39;
    reg PHASE_13;
    wire [63:0] _1167;
    wire [11:0] address_59;
    wire write_enable_59;
    wire [11:0] address_60;
    wire _1354;
    wire read_enable_49;
    wire _1352;
    wire write_enable_60;
    wire _1356;
    wire [131:0] _1361;
    wire [63:0] _1362;
    wire [11:0] _1347 = 12'b000000000000;
    wire [11:0] address_61;
    wire _1345;
    wire write_enable_61;
    wire [63:0] _1270;
    wire [63:0] _1269;
    wire [63:0] _1271;
    wire [63:0] _1267;
    wire [63:0] _1266;
    wire [63:0] q1_4;
    wire [63:0] _1272;
    wire [11:0] address_62;
    wire write_enable_62 = 1'b0;
    wire _1257;
    wire read_enable_50;
    wire [11:0] address_63;
    wire _1253;
    wire read_enable_51;
    wire _1251;
    wire write_enable_63;
    wire _1255;
    wire [131:0] _1262;
    wire [63:0] _1263;
    wire [63:0] data_59 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_60;
    wire [11:0] _1245 = 12'b000000000000;
    wire _1243;
    wire _1242;
    wire _1241;
    wire _1240;
    wire _1239;
    wire _1238;
    wire _1237;
    wire _1236;
    wire _1235;
    wire _1234;
    wire _1233;
    wire _1232;
    wire [11:0] _1244;
    wire [11:0] address_64;
    wire write_enable_64 = 1'b0;
    wire _1229;
    wire read_enable_52;
    wire [63:0] data_61;
    wire [63:0] data_62;
    wire _1226;
    wire _1225;
    wire _1224;
    wire _1223;
    wire _1222;
    wire _1221;
    wire _1220;
    wire _1219;
    wire _1218;
    wire _1217;
    wire _1216;
    wire _1215;
    wire [11:0] _1227;
    wire [11:0] address_65;
    wire _1212;
    wire read_enable_53;
    wire _1210;
    wire write_enable_65;
    wire _1214;
    wire [131:0] _1249;
    wire [63:0] _1250;
    wire _1169 = 1'b0;
    wire _1168 = 1'b0;
    wire _1171;
    wire _43;
    reg PHASE_14;
    wire [63:0] _1264;
    wire [11:0] address_66;
    wire _1202;
    wire read_enable_54;
    wire write_enable_66;
    wire _1204;
    wire [11:0] address_67;
    wire _1197;
    wire read_enable_55;
    wire _1195;
    wire write_enable_67;
    wire _1199;
    wire [131:0] _1207;
    wire [63:0] _1208;
    wire [63:0] _1275;
    wire [63:0] data_63;
    wire [63:0] data_64;
    wire [63:0] data_65;
    wire [63:0] data_66;
    wire [11:0] address_68;
    wire _1188;
    wire read_enable_56;
    wire _1185;
    wire _1186;
    wire write_enable_68;
    wire _1190;
    wire [11:0] address_69;
    wire _1181;
    wire read_enable_57;
    wire _1178;
    wire _1179;
    wire write_enable_69;
    wire _1183;
    wire [131:0] _1193;
    wire [63:0] _1194;
    wire _1176 = 1'b0;
    wire _1175 = 1'b0;
    wire _1276;
    wire _45;
    reg PHASE_15;
    wire [63:0] q0_4;
    wire _1173 = 1'b0;
    wire _1172 = 1'b0;
    reg _1174;
    wire [63:0] _1265;
    wire [191:0] _1274;
    wire [63:0] _1277;
    wire [63:0] data_67;
    wire [63:0] data_68;
    wire [63:0] data_69;
    wire [63:0] data_70;
    wire [11:0] address_70;
    wire _1341;
    wire _1340;
    wire read_enable_58;
    wire _1334 = 1'b0;
    wire _1333 = 1'b0;
    wire _1331 = 1'b0;
    wire _1330 = 1'b0;
    wire _1328 = 1'b0;
    wire _1327 = 1'b0;
    wire _1325 = 1'b0;
    wire _1324 = 1'b0;
    wire _1322 = 1'b0;
    wire _1321 = 1'b0;
    wire _1319 = 1'b0;
    wire _1318 = 1'b0;
    wire _1316 = 1'b0;
    wire _1315 = 1'b0;
    wire _1313 = 1'b0;
    wire _1312 = 1'b0;
    wire _1310 = 1'b0;
    wire _1309 = 1'b0;
    reg _1311;
    reg _1314;
    reg _1317;
    reg _1320;
    reg _1323;
    reg _1326;
    reg _1329;
    reg _1332;
    reg _1335;
    wire _1336;
    wire _1307 = 1'b0;
    wire _1306 = 1'b0;
    wire _1304 = 1'b0;
    wire _1303 = 1'b0;
    wire _1301 = 1'b0;
    wire _1300 = 1'b0;
    wire _1298 = 1'b0;
    wire _1297 = 1'b0;
    wire _1295 = 1'b0;
    wire _1294 = 1'b0;
    wire _1292 = 1'b0;
    wire _1291 = 1'b0;
    wire _1289 = 1'b0;
    wire _1288 = 1'b0;
    wire _1286 = 1'b0;
    wire _1285 = 1'b0;
    wire _1283 = 1'b0;
    wire _1282 = 1'b0;
    reg _1284;
    reg _1287;
    reg _1290;
    reg _1293;
    reg _1296;
    reg _1299;
    reg _1302;
    reg _1305;
    reg _1308;
    wire _1337;
    wire _1338;
    wire write_enable_70;
    wire _1343;
    wire [131:0] _1350;
    wire [63:0] _1351;
    wire _1279 = 1'b0;
    wire _1278 = 1'b0;
    wire _1281;
    wire _47;
    reg PHASE_16;
    wire [63:0] _1363;
    wire [11:0] address_71;
    wire write_enable_71;
    wire [11:0] address_72;
    wire _1550;
    wire read_enable_59;
    wire _1548;
    wire write_enable_72;
    wire _1552;
    wire [131:0] _1557;
    wire [63:0] _1558;
    wire [11:0] _1543 = 12'b000000000000;
    wire [11:0] address_73;
    wire _1541;
    wire write_enable_73;
    wire [63:0] _1466;
    wire [63:0] _1465;
    wire [63:0] _1467;
    wire [63:0] _1463;
    wire [63:0] _1462;
    wire [63:0] q1_5;
    wire [63:0] _1468;
    wire [11:0] address_74;
    wire write_enable_74 = 1'b0;
    wire _1453;
    wire read_enable_60;
    wire [11:0] address_75;
    wire _1449;
    wire read_enable_61;
    wire _1447;
    wire write_enable_75;
    wire _1451;
    wire [131:0] _1458;
    wire [63:0] _1459;
    wire [63:0] data_71 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_72;
    wire [11:0] _1441 = 12'b000000000000;
    wire _1439;
    wire _1438;
    wire _1437;
    wire _1436;
    wire _1435;
    wire _1434;
    wire _1433;
    wire _1432;
    wire _1431;
    wire _1430;
    wire _1429;
    wire _1428;
    wire [11:0] _1440;
    wire [11:0] address_76;
    wire write_enable_76 = 1'b0;
    wire _1425;
    wire read_enable_62;
    wire [63:0] data_73;
    wire [63:0] data_74;
    wire _1422;
    wire _1421;
    wire _1420;
    wire _1419;
    wire _1418;
    wire _1417;
    wire _1416;
    wire _1415;
    wire _1414;
    wire _1413;
    wire _1412;
    wire _1411;
    wire [11:0] _1423;
    wire [11:0] address_77;
    wire _1408;
    wire read_enable_63;
    wire _1406;
    wire write_enable_77;
    wire _1410;
    wire [131:0] _1445;
    wire [63:0] _1446;
    wire _1365 = 1'b0;
    wire _1364 = 1'b0;
    wire _1367;
    wire _51;
    reg PHASE_17;
    wire [63:0] _1460;
    wire [11:0] address_78;
    wire _1398;
    wire read_enable_64;
    wire write_enable_78;
    wire _1400;
    wire [11:0] address_79;
    wire _1393;
    wire read_enable_65;
    wire _1391;
    wire write_enable_79;
    wire _1395;
    wire [131:0] _1403;
    wire [63:0] _1404;
    wire [63:0] _1471;
    wire [63:0] data_75;
    wire [63:0] data_76;
    wire [63:0] data_77;
    wire [63:0] data_78;
    wire [11:0] address_80;
    wire _1384;
    wire read_enable_66;
    wire _1381;
    wire _1382;
    wire write_enable_80;
    wire _1386;
    wire [11:0] address_81;
    wire _1377;
    wire read_enable_67;
    wire _1374;
    wire _1375;
    wire write_enable_81;
    wire _1379;
    wire [131:0] _1389;
    wire [63:0] _1390;
    wire _1372 = 1'b0;
    wire _1371 = 1'b0;
    wire _1472;
    wire _53;
    reg PHASE_18;
    wire [63:0] q0_5;
    wire _1369 = 1'b0;
    wire _1368 = 1'b0;
    reg _1370;
    wire [63:0] _1461;
    wire [191:0] _1470;
    wire [63:0] _1473;
    wire [63:0] data_79;
    wire [63:0] data_80;
    wire [63:0] data_81;
    wire [63:0] data_82;
    wire [11:0] address_82;
    wire _1537;
    wire _1536;
    wire read_enable_68;
    wire _1530 = 1'b0;
    wire _1529 = 1'b0;
    wire _1527 = 1'b0;
    wire _1526 = 1'b0;
    wire _1524 = 1'b0;
    wire _1523 = 1'b0;
    wire _1521 = 1'b0;
    wire _1520 = 1'b0;
    wire _1518 = 1'b0;
    wire _1517 = 1'b0;
    wire _1515 = 1'b0;
    wire _1514 = 1'b0;
    wire _1512 = 1'b0;
    wire _1511 = 1'b0;
    wire _1509 = 1'b0;
    wire _1508 = 1'b0;
    wire _1506 = 1'b0;
    wire _1505 = 1'b0;
    reg _1507;
    reg _1510;
    reg _1513;
    reg _1516;
    reg _1519;
    reg _1522;
    reg _1525;
    reg _1528;
    reg _1531;
    wire _1532;
    wire _1503 = 1'b0;
    wire _1502 = 1'b0;
    wire _1500 = 1'b0;
    wire _1499 = 1'b0;
    wire _1497 = 1'b0;
    wire _1496 = 1'b0;
    wire _1494 = 1'b0;
    wire _1493 = 1'b0;
    wire _1491 = 1'b0;
    wire _1490 = 1'b0;
    wire _1488 = 1'b0;
    wire _1487 = 1'b0;
    wire _1485 = 1'b0;
    wire _1484 = 1'b0;
    wire _1482 = 1'b0;
    wire _1481 = 1'b0;
    wire _1479 = 1'b0;
    wire _1478 = 1'b0;
    reg _1480;
    reg _1483;
    reg _1486;
    reg _1489;
    reg _1492;
    reg _1495;
    reg _1498;
    reg _1501;
    reg _1504;
    wire _1533;
    wire _1534;
    wire write_enable_82;
    wire _1539;
    wire [131:0] _1546;
    wire [63:0] _1547;
    wire _1475 = 1'b0;
    wire _1474 = 1'b0;
    wire _1477;
    wire _55;
    reg PHASE_19;
    wire [63:0] _1559;
    wire [11:0] address_83;
    wire write_enable_83;
    wire [11:0] address_84;
    wire _1746;
    wire read_enable_69;
    wire _1744;
    wire write_enable_84;
    wire _1748;
    wire [131:0] _1753;
    wire [63:0] _1754;
    wire [11:0] _1739 = 12'b000000000000;
    wire [11:0] address_85;
    wire _1737;
    wire write_enable_85;
    wire [3:0] _292;
    wire _291;
    wire _289;
    wire [63:0] _288;
    wire [63:0] _287;
    wire [63:0] _286;
    wire [63:0] _285;
    wire [63:0] _284;
    wire [63:0] _283;
    wire [63:0] _282;
    wire [63:0] _1662;
    wire [63:0] _1661;
    wire [63:0] _1663;
    wire [63:0] _1659;
    wire [63:0] _1658;
    wire [63:0] q1_6;
    wire [63:0] _1664;
    wire [11:0] address_86;
    wire write_enable_86 = 1'b0;
    wire _1649;
    wire read_enable_70;
    wire [11:0] address_87;
    wire _1645;
    wire read_enable_71;
    wire _1643;
    wire write_enable_87;
    wire _1647;
    wire [131:0] _1654;
    wire [63:0] _1655;
    wire [63:0] data_83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_84;
    wire [11:0] _1637 = 12'b000000000000;
    wire _1635;
    wire _1634;
    wire _1633;
    wire _1632;
    wire _1631;
    wire _1630;
    wire _1629;
    wire _1628;
    wire _1627;
    wire _1626;
    wire _1625;
    wire _1624;
    wire [11:0] _1636;
    wire [11:0] address_88;
    wire write_enable_88 = 1'b0;
    wire _1621;
    wire read_enable_72;
    wire [63:0] data_85;
    wire [63:0] data_86;
    wire [11:0] _60;
    wire _1618;
    wire _1617;
    wire _1616;
    wire _1615;
    wire _1614;
    wire _1613;
    wire _1612;
    wire _1611;
    wire _1610;
    wire _1609;
    wire _1608;
    wire _1607;
    wire [11:0] _1619;
    wire [11:0] address_89;
    wire _1604;
    wire read_enable_73;
    wire [7:0] _62;
    wire _1602;
    wire write_enable_89;
    wire _1606;
    wire [131:0] _1641;
    wire [63:0] _1642;
    wire _1561 = 1'b0;
    wire _1560 = 1'b0;
    wire _1563;
    wire _63;
    reg PHASE_20;
    wire [63:0] _1656;
    wire [11:0] address_90;
    wire _1594;
    wire read_enable_74;
    wire write_enable_90;
    wire _1596;
    wire [11:0] address_91;
    wire _1589;
    wire read_enable_75;
    wire _1587;
    wire write_enable_91;
    wire _1591;
    wire [131:0] _1599;
    wire [63:0] _1600;
    wire [63:0] _1667;
    wire [63:0] data_87;
    wire [63:0] data_88;
    wire [63:0] data_89;
    wire [63:0] data_90;
    wire [11:0] _198 = 12'b000000000000;
    wire [11:0] _197 = 12'b000000000000;
    wire [11:0] _195 = 12'b000000000000;
    wire [11:0] _194 = 12'b000000000000;
    wire [11:0] _192 = 12'b000000000000;
    wire [11:0] _191 = 12'b000000000000;
    wire [11:0] _189 = 12'b000000000000;
    wire [11:0] _188 = 12'b000000000000;
    wire [11:0] _186 = 12'b000000000000;
    wire [11:0] _185 = 12'b000000000000;
    wire [11:0] _183 = 12'b000000000000;
    wire [11:0] _182 = 12'b000000000000;
    wire [11:0] _180 = 12'b000000000000;
    wire [11:0] _179 = 12'b000000000000;
    wire [11:0] _177 = 12'b000000000000;
    wire [11:0] _176 = 12'b000000000000;
    wire [11:0] _174 = 12'b000000000000;
    wire [11:0] _173 = 12'b000000000000;
    reg [11:0] _175;
    reg [11:0] _178;
    reg [11:0] _181;
    reg [11:0] _184;
    reg [11:0] _187;
    reg [11:0] _190;
    reg [11:0] _193;
    reg [11:0] _196;
    reg [11:0] _199;
    wire [11:0] _172;
    wire [11:0] address_92;
    wire _1580;
    wire read_enable_76;
    wire _1577;
    wire _1578;
    wire write_enable_92;
    wire _1582;
    wire [11:0] address_93;
    wire _1573;
    wire read_enable_77;
    wire _1570;
    wire _1571;
    wire write_enable_93;
    wire _1575;
    wire [131:0] _1585;
    wire [63:0] _1586;
    wire _99;
    wire _1568 = 1'b0;
    wire _1567 = 1'b0;
    wire _1668;
    wire _65;
    reg PHASE_21;
    wire [63:0] q0_6;
    wire _1565 = 1'b0;
    wire _1564 = 1'b0;
    wire _92;
    reg _1566;
    wire [63:0] _1657;
    wire [191:0] _1666;
    wire [63:0] _1669;
    wire [63:0] data_91;
    wire [63:0] data_92;
    wire [63:0] data_93;
    wire [63:0] data_94;
    wire [11:0] _163 = 12'b000000000000;
    wire [11:0] _162 = 12'b000000000000;
    wire [11:0] _160 = 12'b000000000000;
    wire [11:0] _159 = 12'b000000000000;
    wire [11:0] _157 = 12'b000000000000;
    wire [11:0] _156 = 12'b000000000000;
    wire [11:0] _154 = 12'b000000000000;
    wire [11:0] _153 = 12'b000000000000;
    wire [11:0] _151 = 12'b000000000000;
    wire [11:0] _150 = 12'b000000000000;
    wire [11:0] _148 = 12'b000000000000;
    wire [11:0] _147 = 12'b000000000000;
    wire [11:0] _145 = 12'b000000000000;
    wire [11:0] _144 = 12'b000000000000;
    wire [11:0] _142 = 12'b000000000000;
    wire [11:0] _141 = 12'b000000000000;
    wire [11:0] _139 = 12'b000000000000;
    wire [11:0] _138 = 12'b000000000000;
    wire [11:0] _137;
    reg [11:0] _140;
    reg [11:0] _143;
    reg [11:0] _146;
    reg [11:0] _149;
    reg [11:0] _152;
    reg [11:0] _155;
    reg [11:0] _158;
    reg [11:0] _161;
    reg [11:0] _164;
    wire [11:0] _68;
    wire [11:0] address_94;
    wire _1733;
    wire [7:0] _70;
    wire _1732;
    wire read_enable_78;
    wire _1726 = 1'b0;
    wire _1725 = 1'b0;
    wire _1723 = 1'b0;
    wire _1722 = 1'b0;
    wire _1720 = 1'b0;
    wire _1719 = 1'b0;
    wire _1717 = 1'b0;
    wire _1716 = 1'b0;
    wire _1714 = 1'b0;
    wire _1713 = 1'b0;
    wire _1711 = 1'b0;
    wire _1710 = 1'b0;
    wire _1708 = 1'b0;
    wire _1707 = 1'b0;
    wire _1705 = 1'b0;
    wire _1704 = 1'b0;
    wire _1702 = 1'b0;
    wire _1701 = 1'b0;
    wire _290;
    reg _1703;
    reg _1706;
    reg _1709;
    reg _1712;
    reg _1715;
    reg _1718;
    reg _1721;
    reg _1724;
    reg _1727;
    wire _1728;
    wire _1699 = 1'b0;
    wire _1698 = 1'b0;
    wire _1696 = 1'b0;
    wire _1695 = 1'b0;
    wire _1693 = 1'b0;
    wire _1692 = 1'b0;
    wire _1690 = 1'b0;
    wire _1689 = 1'b0;
    wire _1687 = 1'b0;
    wire _1686 = 1'b0;
    wire _1684 = 1'b0;
    wire _1683 = 1'b0;
    wire _1681 = 1'b0;
    wire _1680 = 1'b0;
    wire _1678 = 1'b0;
    wire _1677 = 1'b0;
    wire _1675 = 1'b0;
    wire _1674 = 1'b0;
    wire _130;
    reg _1676;
    reg _1679;
    reg _1682;
    reg _1685;
    reg _1688;
    reg _1691;
    reg _1694;
    reg _1697;
    reg _1700;
    wire _1729;
    wire _128 = 1'b0;
    wire _127 = 1'b0;
    wire _125 = 1'b0;
    wire _124 = 1'b0;
    wire _122 = 1'b0;
    wire _121 = 1'b0;
    wire _119 = 1'b0;
    wire _118 = 1'b0;
    wire _116 = 1'b0;
    wire _115 = 1'b0;
    wire _113 = 1'b0;
    wire _112 = 1'b0;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire vdd = 1'b1;
    wire _104 = 1'b0;
    wire _103 = 1'b0;
    wire _102;
    reg _105;
    reg _108;
    reg _111;
    reg _114;
    reg _117;
    reg _120;
    reg _123;
    reg _126;
    reg _129;
    wire _1730;
    wire write_enable_94;
    wire _1735;
    wire gnd = 1'b0;
    wire [131:0] _1742;
    wire [63:0] _1743;
    wire _72;
    wire _1671 = 1'b0;
    wire _1670 = 1'b0;
    wire _1673;
    wire _73;
    reg PHASE_22;
    wire [63:0] _1755;
    wire _76;
    wire _78;
    wire _80;
    wire _82;
    wire _84;
    wire [523:0] _91;
    wire _1756;

    /* logic */
    assign address = _372 ? _199 : _367;
    assign write_enable = _365 & _372;
    assign address_0 = _372 ? _164 : _68;
    assign _374 = ~ _372;
    assign read_enable = _360 & _374;
    assign _372 = ~ PHASE_1;
    assign write_enable_0 = _358 & _372;
    assign _376 = write_enable_0 | read_enable;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_376), .regcea(vdd), .wea(write_enable_0), .addra(address_0), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable), .regceb(vdd), .web(write_enable), .addrb(address), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_381[131:131]), .sbiterrb(_381[130:130]), .doutb(_381[129:66]), .dbiterra(_381[65:65]), .sbiterra(_381[64:64]), .douta(_381[63:0]) );
    assign _382 = _381[63:0];
    assign address_1 = PHASE_1 ? _199 : _367;
    assign _365 = _129 & _328;
    assign write_enable_1 = _365 & PHASE_1;
    assign _279 = _271[129:66];
    assign _278 = _258[129:66];
    assign _280 = PHASE ? _279 : _278;
    assign _276 = _216[129:66];
    assign _275 = _202[129:66];
    assign q1 = PHASE_0 ? _276 : _275;
    assign _281 = _96 ? _280 : q1;
    assign address_2 = _260 ? _254 : _253;
    assign _266 = ~ _260;
    assign read_enable_0 = _102 & _266;
    assign address_3 = _260 ? _60 : _236;
    assign _262 = ~ _260;
    assign read_enable_1 = _102 & _262;
    assign _260 = ~ PHASE;
    assign write_enable_3 = _219 & _260;
    assign _264 = write_enable_3 | read_enable_1;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_0
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_264), .regcea(vdd), .wea(write_enable_3), .addra(address_3), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_0), .regceb(vdd), .web(write_enable_2), .addrb(address_2), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_271[131:131]), .sbiterrb(_271[130:130]), .doutb(_271[129:66]), .dbiterra(_271[65:65]), .sbiterra(_271[64:64]), .douta(_271[63:0]) );
    assign _272 = _271[63:0];
    assign _252 = _172[11:11];
    assign _251 = _172[10:10];
    assign _250 = _172[9:9];
    assign _249 = _172[8:8];
    assign _248 = _172[7:7];
    assign _247 = _172[6:6];
    assign _246 = _172[5:5];
    assign _245 = _172[4:4];
    assign _244 = _172[3:3];
    assign _243 = _172[2:2];
    assign _242 = _172[1:1];
    assign _241 = _172[0:0];
    assign _253 = { _241, _242, _243, _244, _245, _246, _247, _248, _249, _250, _251, _252 };
    assign address_4 = PHASE ? _254 : _253;
    assign _238 = ~ PHASE;
    assign read_enable_2 = _102 & _238;
    assign data_1 = wr_d7;
    assign _235 = _137[11:11];
    assign _234 = _137[10:10];
    assign _233 = _137[9:9];
    assign _232 = _137[8:8];
    assign _231 = _137[7:7];
    assign _230 = _137[6:6];
    assign _229 = _137[5:5];
    assign _228 = _137[4:4];
    assign _227 = _137[3:3];
    assign _226 = _137[2:2];
    assign _225 = _137[1:1];
    assign _224 = _137[0:0];
    assign _236 = { _224, _225, _226, _227, _228, _229, _230, _231, _232, _233, _234, _235 };
    assign address_5 = PHASE ? _60 : _236;
    assign _221 = ~ PHASE;
    assign read_enable_3 = _102 & _221;
    assign _219 = _62[7:7];
    assign write_enable_5 = _219 & PHASE;
    assign _223 = write_enable_5 | read_enable_3;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_1
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_223), .regcea(vdd), .wea(write_enable_5), .addra(address_5), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_2), .regceb(vdd), .web(write_enable_4), .addrb(address_4), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_258[131:131]), .sbiterrb(_258[130:130]), .doutb(_258[129:66]), .dbiterra(_258[65:65]), .sbiterra(_258[64:64]), .douta(_258[63:0]) );
    assign _259 = _258[63:0];
    assign _89 = ~ PHASE;
    assign _3 = _89;
    always @(posedge _84) begin
        if (_82)
            PHASE <= _87;
        else
            if (_72)
                PHASE <= _3;
    end
    assign _273 = PHASE ? _272 : _259;
    assign address_6 = _204 ? _199 : _172;
    assign _211 = ~ _204;
    assign read_enable_4 = _102 & _211;
    assign write_enable_6 = _167 & _204;
    assign _213 = write_enable_6 | read_enable_4;
    assign address_7 = _204 ? _164 : _137;
    assign _206 = ~ _204;
    assign read_enable_5 = _102 & _206;
    assign _204 = ~ PHASE_0;
    assign write_enable_7 = _132 & _204;
    assign _208 = write_enable_7 | read_enable_5;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_2
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_208), .regcea(vdd), .wea(write_enable_7), .addra(address_7), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_213), .regceb(vdd), .web(write_enable_6), .addrb(address_6), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_216[131:131]), .sbiterrb(_216[130:130]), .doutb(_216[129:66]), .dbiterra(_216[65:65]), .sbiterra(_216[64:64]), .douta(_216[63:0]) );
    assign _217 = _216[63:0];
    assign _295 = _294[127:64];
    assign data_3 = _295;
    assign address_8 = PHASE_0 ? _199 : _172;
    assign _169 = ~ PHASE_0;
    assign read_enable_6 = _102 & _169;
    assign _166 = ~ _130;
    assign _167 = _129 & _166;
    assign write_enable_8 = _167 & PHASE_0;
    assign _171 = write_enable_8 | read_enable_6;
    assign address_9 = PHASE_0 ? _164 : _137;
    assign _134 = ~ PHASE_0;
    assign read_enable_7 = _102 & _134;
    assign _131 = ~ _130;
    assign _132 = _129 & _131;
    assign write_enable_9 = _132 & PHASE_0;
    assign _136 = write_enable_9 | read_enable_7;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_3
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_136), .regcea(vdd), .wea(write_enable_9), .addra(address_9), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_171), .regceb(vdd), .web(write_enable_8), .addrb(address_8), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_202[131:131]), .sbiterrb(_202[130:130]), .doutb(_202[129:66]), .dbiterra(_202[65:65]), .sbiterra(_202[64:64]), .douta(_202[63:0]) );
    assign _203 = _202[63:0];
    assign _296 = ~ PHASE_0;
    assign _5 = _296;
    always @(posedge _84) begin
        if (_82)
            PHASE_0 <= _98;
        else
            if (_99)
                PHASE_0 <= _5;
    end
    assign q0 = PHASE_0 ? _217 : _203;
    always @(posedge _84) begin
        if (_82)
            _96 <= _94;
        else
            _96 <= _92;
    end
    assign _274 = _96 ? _273 : q0;
    dp_14
        dp_6
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_274), .d2(_281), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_294[191:128]), .q2(_294[127:64]), .q1(_294[63:0]) );
    assign _297 = _294[63:0];
    assign data_7 = _297;
    assign address_10 = PHASE_1 ? _164 : _68;
    assign _361 = ~ PHASE_1;
    assign _360 = _70[7:7];
    assign read_enable_8 = _360 & _361;
    always @(posedge _84) begin
        if (_82)
            _331 <= _330;
        else
            _331 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _334 <= _333;
        else
            _334 <= _331;
    end
    always @(posedge _84) begin
        if (_82)
            _337 <= _336;
        else
            _337 <= _334;
    end
    always @(posedge _84) begin
        if (_82)
            _340 <= _339;
        else
            _340 <= _337;
    end
    always @(posedge _84) begin
        if (_82)
            _343 <= _342;
        else
            _343 <= _340;
    end
    always @(posedge _84) begin
        if (_82)
            _346 <= _345;
        else
            _346 <= _343;
    end
    always @(posedge _84) begin
        if (_82)
            _349 <= _348;
        else
            _349 <= _346;
    end
    always @(posedge _84) begin
        if (_82)
            _352 <= _351;
        else
            _352 <= _349;
    end
    always @(posedge _84) begin
        if (_82)
            _355 <= _354;
        else
            _355 <= _352;
    end
    assign _356 = ~ _355;
    always @(posedge _84) begin
        if (_82)
            _304 <= _303;
        else
            _304 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _307 <= _306;
        else
            _307 <= _304;
    end
    always @(posedge _84) begin
        if (_82)
            _310 <= _309;
        else
            _310 <= _307;
    end
    always @(posedge _84) begin
        if (_82)
            _313 <= _312;
        else
            _313 <= _310;
    end
    always @(posedge _84) begin
        if (_82)
            _316 <= _315;
        else
            _316 <= _313;
    end
    always @(posedge _84) begin
        if (_82)
            _319 <= _318;
        else
            _319 <= _316;
    end
    always @(posedge _84) begin
        if (_82)
            _322 <= _321;
        else
            _322 <= _319;
    end
    always @(posedge _84) begin
        if (_82)
            _325 <= _324;
        else
            _325 <= _322;
    end
    always @(posedge _84) begin
        if (_82)
            _328 <= _327;
        else
            _328 <= _325;
    end
    assign _357 = _328 & _356;
    assign _358 = _129 & _357;
    assign write_enable_10 = _358 & PHASE_1;
    assign _363 = write_enable_10 | read_enable_8;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_4
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_363), .regcea(vdd), .wea(write_enable_10), .addra(address_10), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_1), .regceb(vdd), .web(write_enable_1), .addrb(address_1), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_370[131:131]), .sbiterrb(_370[130:130]), .doutb(_370[129:66]), .dbiterra(_370[65:65]), .sbiterra(_370[64:64]), .douta(_370[63:0]) );
    assign _371 = _370[63:0];
    assign _301 = ~ PHASE_1;
    assign _7 = _301;
    always @(posedge _84) begin
        if (_82)
            PHASE_1 <= _299;
        else
            if (_72)
                PHASE_1 <= _7;
    end
    assign _383 = PHASE_1 ? _382 : _371;
    assign address_11 = _568 ? _199 : _563;
    assign write_enable_11 = _561 & _568;
    assign address_12 = _568 ? _164 : _68;
    assign _570 = ~ _568;
    assign read_enable_9 = _556 & _570;
    assign _568 = ~ PHASE_4;
    assign write_enable_12 = _554 & _568;
    assign _572 = write_enable_12 | read_enable_9;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_5
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_572), .regcea(vdd), .wea(write_enable_12), .addra(address_12), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_11), .regceb(vdd), .web(write_enable_11), .addrb(address_11), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_577[131:131]), .sbiterrb(_577[130:130]), .doutb(_577[129:66]), .dbiterra(_577[65:65]), .sbiterra(_577[64:64]), .douta(_577[63:0]) );
    assign _578 = _577[63:0];
    assign address_13 = PHASE_4 ? _199 : _563;
    assign _561 = _129 & _524;
    assign write_enable_13 = _561 & PHASE_4;
    assign _486 = _478[129:66];
    assign _485 = _465[129:66];
    assign _487 = PHASE_2 ? _486 : _485;
    assign _483 = _423[129:66];
    assign _482 = _409[129:66];
    assign q1_0 = PHASE_3 ? _483 : _482;
    assign _488 = _390 ? _487 : q1_0;
    assign address_14 = _467 ? _461 : _460;
    assign _473 = ~ _467;
    assign read_enable_10 = _102 & _473;
    assign address_15 = _467 ? _60 : _443;
    assign _469 = ~ _467;
    assign read_enable_11 = _102 & _469;
    assign _467 = ~ PHASE_2;
    assign write_enable_15 = _426 & _467;
    assign _471 = write_enable_15 | read_enable_11;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_6
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_471), .regcea(vdd), .wea(write_enable_15), .addra(address_15), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_10), .regceb(vdd), .web(write_enable_14), .addrb(address_14), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_478[131:131]), .sbiterrb(_478[130:130]), .doutb(_478[129:66]), .dbiterra(_478[65:65]), .sbiterra(_478[64:64]), .douta(_478[63:0]) );
    assign _479 = _478[63:0];
    assign _459 = _172[11:11];
    assign _458 = _172[10:10];
    assign _457 = _172[9:9];
    assign _456 = _172[8:8];
    assign _455 = _172[7:7];
    assign _454 = _172[6:6];
    assign _453 = _172[5:5];
    assign _452 = _172[4:4];
    assign _451 = _172[3:3];
    assign _450 = _172[2:2];
    assign _449 = _172[1:1];
    assign _448 = _172[0:0];
    assign _460 = { _448, _449, _450, _451, _452, _453, _454, _455, _456, _457, _458, _459 };
    assign address_16 = PHASE_2 ? _461 : _460;
    assign _445 = ~ PHASE_2;
    assign read_enable_12 = _102 & _445;
    assign data_13 = wr_d6;
    assign _442 = _137[11:11];
    assign _441 = _137[10:10];
    assign _440 = _137[9:9];
    assign _439 = _137[8:8];
    assign _438 = _137[7:7];
    assign _437 = _137[6:6];
    assign _436 = _137[5:5];
    assign _435 = _137[4:4];
    assign _434 = _137[3:3];
    assign _433 = _137[2:2];
    assign _432 = _137[1:1];
    assign _431 = _137[0:0];
    assign _443 = { _431, _432, _433, _434, _435, _436, _437, _438, _439, _440, _441, _442 };
    assign address_17 = PHASE_2 ? _60 : _443;
    assign _428 = ~ PHASE_2;
    assign read_enable_13 = _102 & _428;
    assign _426 = _62[6:6];
    assign write_enable_17 = _426 & PHASE_2;
    assign _430 = write_enable_17 | read_enable_13;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_7
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_430), .regcea(vdd), .wea(write_enable_17), .addra(address_17), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_12), .regceb(vdd), .web(write_enable_16), .addrb(address_16), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_465[131:131]), .sbiterrb(_465[130:130]), .doutb(_465[129:66]), .dbiterra(_465[65:65]), .sbiterra(_465[64:64]), .douta(_465[63:0]) );
    assign _466 = _465[63:0];
    assign _387 = ~ PHASE_2;
    assign _11 = _387;
    always @(posedge _84) begin
        if (_82)
            PHASE_2 <= _385;
        else
            if (_72)
                PHASE_2 <= _11;
    end
    assign _480 = PHASE_2 ? _479 : _466;
    assign address_18 = _411 ? _199 : _172;
    assign _418 = ~ _411;
    assign read_enable_14 = _102 & _418;
    assign write_enable_18 = _402 & _411;
    assign _420 = write_enable_18 | read_enable_14;
    assign address_19 = _411 ? _164 : _137;
    assign _413 = ~ _411;
    assign read_enable_15 = _102 & _413;
    assign _411 = ~ PHASE_3;
    assign write_enable_19 = _395 & _411;
    assign _415 = write_enable_19 | read_enable_15;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_8
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_415), .regcea(vdd), .wea(write_enable_19), .addra(address_19), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_420), .regceb(vdd), .web(write_enable_18), .addrb(address_18), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_423[131:131]), .sbiterrb(_423[130:130]), .doutb(_423[129:66]), .dbiterra(_423[65:65]), .sbiterra(_423[64:64]), .douta(_423[63:0]) );
    assign _424 = _423[63:0];
    assign _491 = _490[127:64];
    assign data_15 = _491;
    assign address_20 = PHASE_3 ? _199 : _172;
    assign _404 = ~ PHASE_3;
    assign read_enable_16 = _102 & _404;
    assign _401 = ~ _130;
    assign _402 = _129 & _401;
    assign write_enable_20 = _402 & PHASE_3;
    assign _406 = write_enable_20 | read_enable_16;
    assign address_21 = PHASE_3 ? _164 : _137;
    assign _397 = ~ PHASE_3;
    assign read_enable_17 = _102 & _397;
    assign _394 = ~ _130;
    assign _395 = _129 & _394;
    assign write_enable_21 = _395 & PHASE_3;
    assign _399 = write_enable_21 | read_enable_17;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_9
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_399), .regcea(vdd), .wea(write_enable_21), .addra(address_21), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_406), .regceb(vdd), .web(write_enable_20), .addrb(address_20), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_409[131:131]), .sbiterrb(_409[130:130]), .doutb(_409[129:66]), .dbiterra(_409[65:65]), .sbiterra(_409[64:64]), .douta(_409[63:0]) );
    assign _410 = _409[63:0];
    assign _492 = ~ PHASE_3;
    assign _13 = _492;
    always @(posedge _84) begin
        if (_82)
            PHASE_3 <= _392;
        else
            if (_99)
                PHASE_3 <= _13;
    end
    assign q0_0 = PHASE_3 ? _424 : _410;
    always @(posedge _84) begin
        if (_82)
            _390 <= _389;
        else
            _390 <= _92;
    end
    assign _481 = _390 ? _480 : q0_0;
    dp_13
        dp_5
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_481), .d2(_488), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_490[191:128]), .q2(_490[127:64]), .q1(_490[63:0]) );
    assign _493 = _490[63:0];
    assign data_19 = _493;
    assign address_22 = PHASE_4 ? _164 : _68;
    assign _557 = ~ PHASE_4;
    assign _556 = _70[6:6];
    assign read_enable_18 = _556 & _557;
    always @(posedge _84) begin
        if (_82)
            _527 <= _526;
        else
            _527 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _530 <= _529;
        else
            _530 <= _527;
    end
    always @(posedge _84) begin
        if (_82)
            _533 <= _532;
        else
            _533 <= _530;
    end
    always @(posedge _84) begin
        if (_82)
            _536 <= _535;
        else
            _536 <= _533;
    end
    always @(posedge _84) begin
        if (_82)
            _539 <= _538;
        else
            _539 <= _536;
    end
    always @(posedge _84) begin
        if (_82)
            _542 <= _541;
        else
            _542 <= _539;
    end
    always @(posedge _84) begin
        if (_82)
            _545 <= _544;
        else
            _545 <= _542;
    end
    always @(posedge _84) begin
        if (_82)
            _548 <= _547;
        else
            _548 <= _545;
    end
    always @(posedge _84) begin
        if (_82)
            _551 <= _550;
        else
            _551 <= _548;
    end
    assign _552 = ~ _551;
    always @(posedge _84) begin
        if (_82)
            _500 <= _499;
        else
            _500 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _503 <= _502;
        else
            _503 <= _500;
    end
    always @(posedge _84) begin
        if (_82)
            _506 <= _505;
        else
            _506 <= _503;
    end
    always @(posedge _84) begin
        if (_82)
            _509 <= _508;
        else
            _509 <= _506;
    end
    always @(posedge _84) begin
        if (_82)
            _512 <= _511;
        else
            _512 <= _509;
    end
    always @(posedge _84) begin
        if (_82)
            _515 <= _514;
        else
            _515 <= _512;
    end
    always @(posedge _84) begin
        if (_82)
            _518 <= _517;
        else
            _518 <= _515;
    end
    always @(posedge _84) begin
        if (_82)
            _521 <= _520;
        else
            _521 <= _518;
    end
    always @(posedge _84) begin
        if (_82)
            _524 <= _523;
        else
            _524 <= _521;
    end
    assign _553 = _524 & _552;
    assign _554 = _129 & _553;
    assign write_enable_22 = _554 & PHASE_4;
    assign _559 = write_enable_22 | read_enable_18;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_10
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_559), .regcea(vdd), .wea(write_enable_22), .addra(address_22), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_13), .regceb(vdd), .web(write_enable_13), .addrb(address_13), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_566[131:131]), .sbiterrb(_566[130:130]), .doutb(_566[129:66]), .dbiterra(_566[65:65]), .sbiterra(_566[64:64]), .douta(_566[63:0]) );
    assign _567 = _566[63:0];
    assign _497 = ~ PHASE_4;
    assign _15 = _497;
    always @(posedge _84) begin
        if (_82)
            PHASE_4 <= _495;
        else
            if (_72)
                PHASE_4 <= _15;
    end
    assign _579 = PHASE_4 ? _578 : _567;
    assign address_23 = _764 ? _199 : _759;
    assign write_enable_23 = _757 & _764;
    assign address_24 = _764 ? _164 : _68;
    assign _766 = ~ _764;
    assign read_enable_19 = _752 & _766;
    assign _764 = ~ PHASE_7;
    assign write_enable_24 = _750 & _764;
    assign _768 = write_enable_24 | read_enable_19;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_11
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_768), .regcea(vdd), .wea(write_enable_24), .addra(address_24), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_23), .regceb(vdd), .web(write_enable_23), .addrb(address_23), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_773[131:131]), .sbiterrb(_773[130:130]), .doutb(_773[129:66]), .dbiterra(_773[65:65]), .sbiterra(_773[64:64]), .douta(_773[63:0]) );
    assign _774 = _773[63:0];
    assign address_25 = PHASE_7 ? _199 : _759;
    assign _757 = _129 & _720;
    assign write_enable_25 = _757 & PHASE_7;
    assign _682 = _674[129:66];
    assign _681 = _661[129:66];
    assign _683 = PHASE_5 ? _682 : _681;
    assign _679 = _619[129:66];
    assign _678 = _605[129:66];
    assign q1_1 = PHASE_6 ? _679 : _678;
    assign _684 = _586 ? _683 : q1_1;
    assign address_26 = _663 ? _657 : _656;
    assign _669 = ~ _663;
    assign read_enable_20 = _102 & _669;
    assign address_27 = _663 ? _60 : _639;
    assign _665 = ~ _663;
    assign read_enable_21 = _102 & _665;
    assign _663 = ~ PHASE_5;
    assign write_enable_27 = _622 & _663;
    assign _667 = write_enable_27 | read_enable_21;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_12
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_667), .regcea(vdd), .wea(write_enable_27), .addra(address_27), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_20), .regceb(vdd), .web(write_enable_26), .addrb(address_26), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_674[131:131]), .sbiterrb(_674[130:130]), .doutb(_674[129:66]), .dbiterra(_674[65:65]), .sbiterra(_674[64:64]), .douta(_674[63:0]) );
    assign _675 = _674[63:0];
    assign _655 = _172[11:11];
    assign _654 = _172[10:10];
    assign _653 = _172[9:9];
    assign _652 = _172[8:8];
    assign _651 = _172[7:7];
    assign _650 = _172[6:6];
    assign _649 = _172[5:5];
    assign _648 = _172[4:4];
    assign _647 = _172[3:3];
    assign _646 = _172[2:2];
    assign _645 = _172[1:1];
    assign _644 = _172[0:0];
    assign _656 = { _644, _645, _646, _647, _648, _649, _650, _651, _652, _653, _654, _655 };
    assign address_28 = PHASE_5 ? _657 : _656;
    assign _641 = ~ PHASE_5;
    assign read_enable_22 = _102 & _641;
    assign data_25 = wr_d5;
    assign _638 = _137[11:11];
    assign _637 = _137[10:10];
    assign _636 = _137[9:9];
    assign _635 = _137[8:8];
    assign _634 = _137[7:7];
    assign _633 = _137[6:6];
    assign _632 = _137[5:5];
    assign _631 = _137[4:4];
    assign _630 = _137[3:3];
    assign _629 = _137[2:2];
    assign _628 = _137[1:1];
    assign _627 = _137[0:0];
    assign _639 = { _627, _628, _629, _630, _631, _632, _633, _634, _635, _636, _637, _638 };
    assign address_29 = PHASE_5 ? _60 : _639;
    assign _624 = ~ PHASE_5;
    assign read_enable_23 = _102 & _624;
    assign _622 = _62[5:5];
    assign write_enable_29 = _622 & PHASE_5;
    assign _626 = write_enable_29 | read_enable_23;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_13
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_626), .regcea(vdd), .wea(write_enable_29), .addra(address_29), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_22), .regceb(vdd), .web(write_enable_28), .addrb(address_28), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_661[131:131]), .sbiterrb(_661[130:130]), .doutb(_661[129:66]), .dbiterra(_661[65:65]), .sbiterra(_661[64:64]), .douta(_661[63:0]) );
    assign _662 = _661[63:0];
    assign _583 = ~ PHASE_5;
    assign _19 = _583;
    always @(posedge _84) begin
        if (_82)
            PHASE_5 <= _581;
        else
            if (_72)
                PHASE_5 <= _19;
    end
    assign _676 = PHASE_5 ? _675 : _662;
    assign address_30 = _607 ? _199 : _172;
    assign _614 = ~ _607;
    assign read_enable_24 = _102 & _614;
    assign write_enable_30 = _598 & _607;
    assign _616 = write_enable_30 | read_enable_24;
    assign address_31 = _607 ? _164 : _137;
    assign _609 = ~ _607;
    assign read_enable_25 = _102 & _609;
    assign _607 = ~ PHASE_6;
    assign write_enable_31 = _591 & _607;
    assign _611 = write_enable_31 | read_enable_25;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_14
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_611), .regcea(vdd), .wea(write_enable_31), .addra(address_31), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_616), .regceb(vdd), .web(write_enable_30), .addrb(address_30), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_619[131:131]), .sbiterrb(_619[130:130]), .doutb(_619[129:66]), .dbiterra(_619[65:65]), .sbiterra(_619[64:64]), .douta(_619[63:0]) );
    assign _620 = _619[63:0];
    assign _687 = _686[127:64];
    assign data_27 = _687;
    assign address_32 = PHASE_6 ? _199 : _172;
    assign _600 = ~ PHASE_6;
    assign read_enable_26 = _102 & _600;
    assign _597 = ~ _130;
    assign _598 = _129 & _597;
    assign write_enable_32 = _598 & PHASE_6;
    assign _602 = write_enable_32 | read_enable_26;
    assign address_33 = PHASE_6 ? _164 : _137;
    assign _593 = ~ PHASE_6;
    assign read_enable_27 = _102 & _593;
    assign _590 = ~ _130;
    assign _591 = _129 & _590;
    assign write_enable_33 = _591 & PHASE_6;
    assign _595 = write_enable_33 | read_enable_27;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_15
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_595), .regcea(vdd), .wea(write_enable_33), .addra(address_33), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_602), .regceb(vdd), .web(write_enable_32), .addrb(address_32), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_605[131:131]), .sbiterrb(_605[130:130]), .doutb(_605[129:66]), .dbiterra(_605[65:65]), .sbiterra(_605[64:64]), .douta(_605[63:0]) );
    assign _606 = _605[63:0];
    assign _688 = ~ PHASE_6;
    assign _21 = _688;
    always @(posedge _84) begin
        if (_82)
            PHASE_6 <= _588;
        else
            if (_99)
                PHASE_6 <= _21;
    end
    assign q0_1 = PHASE_6 ? _620 : _606;
    always @(posedge _84) begin
        if (_82)
            _586 <= _585;
        else
            _586 <= _92;
    end
    assign _677 = _586 ? _676 : q0_1;
    dp_12
        dp_4
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_677), .d2(_684), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_686[191:128]), .q2(_686[127:64]), .q1(_686[63:0]) );
    assign _689 = _686[63:0];
    assign data_31 = _689;
    assign address_34 = PHASE_7 ? _164 : _68;
    assign _753 = ~ PHASE_7;
    assign _752 = _70[5:5];
    assign read_enable_28 = _752 & _753;
    always @(posedge _84) begin
        if (_82)
            _723 <= _722;
        else
            _723 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _726 <= _725;
        else
            _726 <= _723;
    end
    always @(posedge _84) begin
        if (_82)
            _729 <= _728;
        else
            _729 <= _726;
    end
    always @(posedge _84) begin
        if (_82)
            _732 <= _731;
        else
            _732 <= _729;
    end
    always @(posedge _84) begin
        if (_82)
            _735 <= _734;
        else
            _735 <= _732;
    end
    always @(posedge _84) begin
        if (_82)
            _738 <= _737;
        else
            _738 <= _735;
    end
    always @(posedge _84) begin
        if (_82)
            _741 <= _740;
        else
            _741 <= _738;
    end
    always @(posedge _84) begin
        if (_82)
            _744 <= _743;
        else
            _744 <= _741;
    end
    always @(posedge _84) begin
        if (_82)
            _747 <= _746;
        else
            _747 <= _744;
    end
    assign _748 = ~ _747;
    always @(posedge _84) begin
        if (_82)
            _696 <= _695;
        else
            _696 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _699 <= _698;
        else
            _699 <= _696;
    end
    always @(posedge _84) begin
        if (_82)
            _702 <= _701;
        else
            _702 <= _699;
    end
    always @(posedge _84) begin
        if (_82)
            _705 <= _704;
        else
            _705 <= _702;
    end
    always @(posedge _84) begin
        if (_82)
            _708 <= _707;
        else
            _708 <= _705;
    end
    always @(posedge _84) begin
        if (_82)
            _711 <= _710;
        else
            _711 <= _708;
    end
    always @(posedge _84) begin
        if (_82)
            _714 <= _713;
        else
            _714 <= _711;
    end
    always @(posedge _84) begin
        if (_82)
            _717 <= _716;
        else
            _717 <= _714;
    end
    always @(posedge _84) begin
        if (_82)
            _720 <= _719;
        else
            _720 <= _717;
    end
    assign _749 = _720 & _748;
    assign _750 = _129 & _749;
    assign write_enable_34 = _750 & PHASE_7;
    assign _755 = write_enable_34 | read_enable_28;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_16
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_755), .regcea(vdd), .wea(write_enable_34), .addra(address_34), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_25), .regceb(vdd), .web(write_enable_25), .addrb(address_25), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_762[131:131]), .sbiterrb(_762[130:130]), .doutb(_762[129:66]), .dbiterra(_762[65:65]), .sbiterra(_762[64:64]), .douta(_762[63:0]) );
    assign _763 = _762[63:0];
    assign _693 = ~ PHASE_7;
    assign _23 = _693;
    always @(posedge _84) begin
        if (_82)
            PHASE_7 <= _691;
        else
            if (_72)
                PHASE_7 <= _23;
    end
    assign _775 = PHASE_7 ? _774 : _763;
    assign address_35 = _960 ? _199 : _955;
    assign write_enable_35 = _953 & _960;
    assign address_36 = _960 ? _164 : _68;
    assign _962 = ~ _960;
    assign read_enable_29 = _948 & _962;
    assign _960 = ~ PHASE_10;
    assign write_enable_36 = _946 & _960;
    assign _964 = write_enable_36 | read_enable_29;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_17
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_964), .regcea(vdd), .wea(write_enable_36), .addra(address_36), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_35), .regceb(vdd), .web(write_enable_35), .addrb(address_35), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_969[131:131]), .sbiterrb(_969[130:130]), .doutb(_969[129:66]), .dbiterra(_969[65:65]), .sbiterra(_969[64:64]), .douta(_969[63:0]) );
    assign _970 = _969[63:0];
    assign address_37 = PHASE_10 ? _199 : _955;
    assign _953 = _129 & _916;
    assign write_enable_37 = _953 & PHASE_10;
    assign _878 = _870[129:66];
    assign _877 = _857[129:66];
    assign _879 = PHASE_8 ? _878 : _877;
    assign _875 = _815[129:66];
    assign _874 = _801[129:66];
    assign q1_2 = PHASE_9 ? _875 : _874;
    assign _880 = _782 ? _879 : q1_2;
    assign address_38 = _859 ? _853 : _852;
    assign _865 = ~ _859;
    assign read_enable_30 = _102 & _865;
    assign address_39 = _859 ? _60 : _835;
    assign _861 = ~ _859;
    assign read_enable_31 = _102 & _861;
    assign _859 = ~ PHASE_8;
    assign write_enable_39 = _818 & _859;
    assign _863 = write_enable_39 | read_enable_31;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_18
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_863), .regcea(vdd), .wea(write_enable_39), .addra(address_39), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_30), .regceb(vdd), .web(write_enable_38), .addrb(address_38), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_870[131:131]), .sbiterrb(_870[130:130]), .doutb(_870[129:66]), .dbiterra(_870[65:65]), .sbiterra(_870[64:64]), .douta(_870[63:0]) );
    assign _871 = _870[63:0];
    assign _851 = _172[11:11];
    assign _850 = _172[10:10];
    assign _849 = _172[9:9];
    assign _848 = _172[8:8];
    assign _847 = _172[7:7];
    assign _846 = _172[6:6];
    assign _845 = _172[5:5];
    assign _844 = _172[4:4];
    assign _843 = _172[3:3];
    assign _842 = _172[2:2];
    assign _841 = _172[1:1];
    assign _840 = _172[0:0];
    assign _852 = { _840, _841, _842, _843, _844, _845, _846, _847, _848, _849, _850, _851 };
    assign address_40 = PHASE_8 ? _853 : _852;
    assign _837 = ~ PHASE_8;
    assign read_enable_32 = _102 & _837;
    assign data_37 = wr_d4;
    assign _834 = _137[11:11];
    assign _833 = _137[10:10];
    assign _832 = _137[9:9];
    assign _831 = _137[8:8];
    assign _830 = _137[7:7];
    assign _829 = _137[6:6];
    assign _828 = _137[5:5];
    assign _827 = _137[4:4];
    assign _826 = _137[3:3];
    assign _825 = _137[2:2];
    assign _824 = _137[1:1];
    assign _823 = _137[0:0];
    assign _835 = { _823, _824, _825, _826, _827, _828, _829, _830, _831, _832, _833, _834 };
    assign address_41 = PHASE_8 ? _60 : _835;
    assign _820 = ~ PHASE_8;
    assign read_enable_33 = _102 & _820;
    assign _818 = _62[4:4];
    assign write_enable_41 = _818 & PHASE_8;
    assign _822 = write_enable_41 | read_enable_33;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_19
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_822), .regcea(vdd), .wea(write_enable_41), .addra(address_41), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_32), .regceb(vdd), .web(write_enable_40), .addrb(address_40), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_857[131:131]), .sbiterrb(_857[130:130]), .doutb(_857[129:66]), .dbiterra(_857[65:65]), .sbiterra(_857[64:64]), .douta(_857[63:0]) );
    assign _858 = _857[63:0];
    assign _779 = ~ PHASE_8;
    assign _27 = _779;
    always @(posedge _84) begin
        if (_82)
            PHASE_8 <= _777;
        else
            if (_72)
                PHASE_8 <= _27;
    end
    assign _872 = PHASE_8 ? _871 : _858;
    assign address_42 = _803 ? _199 : _172;
    assign _810 = ~ _803;
    assign read_enable_34 = _102 & _810;
    assign write_enable_42 = _794 & _803;
    assign _812 = write_enable_42 | read_enable_34;
    assign address_43 = _803 ? _164 : _137;
    assign _805 = ~ _803;
    assign read_enable_35 = _102 & _805;
    assign _803 = ~ PHASE_9;
    assign write_enable_43 = _787 & _803;
    assign _807 = write_enable_43 | read_enable_35;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_20
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_807), .regcea(vdd), .wea(write_enable_43), .addra(address_43), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_812), .regceb(vdd), .web(write_enable_42), .addrb(address_42), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_815[131:131]), .sbiterrb(_815[130:130]), .doutb(_815[129:66]), .dbiterra(_815[65:65]), .sbiterra(_815[64:64]), .douta(_815[63:0]) );
    assign _816 = _815[63:0];
    assign _883 = _882[127:64];
    assign data_39 = _883;
    assign address_44 = PHASE_9 ? _199 : _172;
    assign _796 = ~ PHASE_9;
    assign read_enable_36 = _102 & _796;
    assign _793 = ~ _130;
    assign _794 = _129 & _793;
    assign write_enable_44 = _794 & PHASE_9;
    assign _798 = write_enable_44 | read_enable_36;
    assign address_45 = PHASE_9 ? _164 : _137;
    assign _789 = ~ PHASE_9;
    assign read_enable_37 = _102 & _789;
    assign _786 = ~ _130;
    assign _787 = _129 & _786;
    assign write_enable_45 = _787 & PHASE_9;
    assign _791 = write_enable_45 | read_enable_37;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_21
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_791), .regcea(vdd), .wea(write_enable_45), .addra(address_45), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_798), .regceb(vdd), .web(write_enable_44), .addrb(address_44), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_801[131:131]), .sbiterrb(_801[130:130]), .doutb(_801[129:66]), .dbiterra(_801[65:65]), .sbiterra(_801[64:64]), .douta(_801[63:0]) );
    assign _802 = _801[63:0];
    assign _884 = ~ PHASE_9;
    assign _29 = _884;
    always @(posedge _84) begin
        if (_82)
            PHASE_9 <= _784;
        else
            if (_99)
                PHASE_9 <= _29;
    end
    assign q0_2 = PHASE_9 ? _816 : _802;
    always @(posedge _84) begin
        if (_82)
            _782 <= _781;
        else
            _782 <= _92;
    end
    assign _873 = _782 ? _872 : q0_2;
    dp_11
        dp_3
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_873), .d2(_880), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_882[191:128]), .q2(_882[127:64]), .q1(_882[63:0]) );
    assign _885 = _882[63:0];
    assign data_43 = _885;
    assign address_46 = PHASE_10 ? _164 : _68;
    assign _949 = ~ PHASE_10;
    assign _948 = _70[4:4];
    assign read_enable_38 = _948 & _949;
    always @(posedge _84) begin
        if (_82)
            _919 <= _918;
        else
            _919 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _922 <= _921;
        else
            _922 <= _919;
    end
    always @(posedge _84) begin
        if (_82)
            _925 <= _924;
        else
            _925 <= _922;
    end
    always @(posedge _84) begin
        if (_82)
            _928 <= _927;
        else
            _928 <= _925;
    end
    always @(posedge _84) begin
        if (_82)
            _931 <= _930;
        else
            _931 <= _928;
    end
    always @(posedge _84) begin
        if (_82)
            _934 <= _933;
        else
            _934 <= _931;
    end
    always @(posedge _84) begin
        if (_82)
            _937 <= _936;
        else
            _937 <= _934;
    end
    always @(posedge _84) begin
        if (_82)
            _940 <= _939;
        else
            _940 <= _937;
    end
    always @(posedge _84) begin
        if (_82)
            _943 <= _942;
        else
            _943 <= _940;
    end
    assign _944 = ~ _943;
    always @(posedge _84) begin
        if (_82)
            _892 <= _891;
        else
            _892 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _895 <= _894;
        else
            _895 <= _892;
    end
    always @(posedge _84) begin
        if (_82)
            _898 <= _897;
        else
            _898 <= _895;
    end
    always @(posedge _84) begin
        if (_82)
            _901 <= _900;
        else
            _901 <= _898;
    end
    always @(posedge _84) begin
        if (_82)
            _904 <= _903;
        else
            _904 <= _901;
    end
    always @(posedge _84) begin
        if (_82)
            _907 <= _906;
        else
            _907 <= _904;
    end
    always @(posedge _84) begin
        if (_82)
            _910 <= _909;
        else
            _910 <= _907;
    end
    always @(posedge _84) begin
        if (_82)
            _913 <= _912;
        else
            _913 <= _910;
    end
    always @(posedge _84) begin
        if (_82)
            _916 <= _915;
        else
            _916 <= _913;
    end
    assign _945 = _916 & _944;
    assign _946 = _129 & _945;
    assign write_enable_46 = _946 & PHASE_10;
    assign _951 = write_enable_46 | read_enable_38;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_22
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_951), .regcea(vdd), .wea(write_enable_46), .addra(address_46), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_37), .regceb(vdd), .web(write_enable_37), .addrb(address_37), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_958[131:131]), .sbiterrb(_958[130:130]), .doutb(_958[129:66]), .dbiterra(_958[65:65]), .sbiterra(_958[64:64]), .douta(_958[63:0]) );
    assign _959 = _958[63:0];
    assign _889 = ~ PHASE_10;
    assign _31 = _889;
    always @(posedge _84) begin
        if (_82)
            PHASE_10 <= _887;
        else
            if (_72)
                PHASE_10 <= _31;
    end
    assign _971 = PHASE_10 ? _970 : _959;
    assign address_47 = _1156 ? _199 : _1151;
    assign write_enable_47 = _1149 & _1156;
    assign address_48 = _1156 ? _164 : _68;
    assign _1158 = ~ _1156;
    assign read_enable_39 = _1144 & _1158;
    assign _1156 = ~ PHASE_13;
    assign write_enable_48 = _1142 & _1156;
    assign _1160 = write_enable_48 | read_enable_39;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_23
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1160), .regcea(vdd), .wea(write_enable_48), .addra(address_48), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_47), .regceb(vdd), .web(write_enable_47), .addrb(address_47), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1165[131:131]), .sbiterrb(_1165[130:130]), .doutb(_1165[129:66]), .dbiterra(_1165[65:65]), .sbiterra(_1165[64:64]), .douta(_1165[63:0]) );
    assign _1166 = _1165[63:0];
    assign address_49 = PHASE_13 ? _199 : _1151;
    assign _1149 = _129 & _1112;
    assign write_enable_49 = _1149 & PHASE_13;
    assign _1074 = _1066[129:66];
    assign _1073 = _1053[129:66];
    assign _1075 = PHASE_11 ? _1074 : _1073;
    assign _1071 = _1011[129:66];
    assign _1070 = _997[129:66];
    assign q1_3 = PHASE_12 ? _1071 : _1070;
    assign _1076 = _978 ? _1075 : q1_3;
    assign address_50 = _1055 ? _1049 : _1048;
    assign _1061 = ~ _1055;
    assign read_enable_40 = _102 & _1061;
    assign address_51 = _1055 ? _60 : _1031;
    assign _1057 = ~ _1055;
    assign read_enable_41 = _102 & _1057;
    assign _1055 = ~ PHASE_11;
    assign write_enable_51 = _1014 & _1055;
    assign _1059 = write_enable_51 | read_enable_41;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_24
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1059), .regcea(vdd), .wea(write_enable_51), .addra(address_51), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_40), .regceb(vdd), .web(write_enable_50), .addrb(address_50), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1066[131:131]), .sbiterrb(_1066[130:130]), .doutb(_1066[129:66]), .dbiterra(_1066[65:65]), .sbiterra(_1066[64:64]), .douta(_1066[63:0]) );
    assign _1067 = _1066[63:0];
    assign _1047 = _172[11:11];
    assign _1046 = _172[10:10];
    assign _1045 = _172[9:9];
    assign _1044 = _172[8:8];
    assign _1043 = _172[7:7];
    assign _1042 = _172[6:6];
    assign _1041 = _172[5:5];
    assign _1040 = _172[4:4];
    assign _1039 = _172[3:3];
    assign _1038 = _172[2:2];
    assign _1037 = _172[1:1];
    assign _1036 = _172[0:0];
    assign _1048 = { _1036, _1037, _1038, _1039, _1040, _1041, _1042, _1043, _1044, _1045, _1046, _1047 };
    assign address_52 = PHASE_11 ? _1049 : _1048;
    assign _1033 = ~ PHASE_11;
    assign read_enable_42 = _102 & _1033;
    assign data_49 = wr_d3;
    assign _1030 = _137[11:11];
    assign _1029 = _137[10:10];
    assign _1028 = _137[9:9];
    assign _1027 = _137[8:8];
    assign _1026 = _137[7:7];
    assign _1025 = _137[6:6];
    assign _1024 = _137[5:5];
    assign _1023 = _137[4:4];
    assign _1022 = _137[3:3];
    assign _1021 = _137[2:2];
    assign _1020 = _137[1:1];
    assign _1019 = _137[0:0];
    assign _1031 = { _1019, _1020, _1021, _1022, _1023, _1024, _1025, _1026, _1027, _1028, _1029, _1030 };
    assign address_53 = PHASE_11 ? _60 : _1031;
    assign _1016 = ~ PHASE_11;
    assign read_enable_43 = _102 & _1016;
    assign _1014 = _62[3:3];
    assign write_enable_53 = _1014 & PHASE_11;
    assign _1018 = write_enable_53 | read_enable_43;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_25
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1018), .regcea(vdd), .wea(write_enable_53), .addra(address_53), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_42), .regceb(vdd), .web(write_enable_52), .addrb(address_52), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1053[131:131]), .sbiterrb(_1053[130:130]), .doutb(_1053[129:66]), .dbiterra(_1053[65:65]), .sbiterra(_1053[64:64]), .douta(_1053[63:0]) );
    assign _1054 = _1053[63:0];
    assign _975 = ~ PHASE_11;
    assign _35 = _975;
    always @(posedge _84) begin
        if (_82)
            PHASE_11 <= _973;
        else
            if (_72)
                PHASE_11 <= _35;
    end
    assign _1068 = PHASE_11 ? _1067 : _1054;
    assign address_54 = _999 ? _199 : _172;
    assign _1006 = ~ _999;
    assign read_enable_44 = _102 & _1006;
    assign write_enable_54 = _990 & _999;
    assign _1008 = write_enable_54 | read_enable_44;
    assign address_55 = _999 ? _164 : _137;
    assign _1001 = ~ _999;
    assign read_enable_45 = _102 & _1001;
    assign _999 = ~ PHASE_12;
    assign write_enable_55 = _983 & _999;
    assign _1003 = write_enable_55 | read_enable_45;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_26
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1003), .regcea(vdd), .wea(write_enable_55), .addra(address_55), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1008), .regceb(vdd), .web(write_enable_54), .addrb(address_54), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1011[131:131]), .sbiterrb(_1011[130:130]), .doutb(_1011[129:66]), .dbiterra(_1011[65:65]), .sbiterra(_1011[64:64]), .douta(_1011[63:0]) );
    assign _1012 = _1011[63:0];
    assign _1079 = _1078[127:64];
    assign data_51 = _1079;
    assign address_56 = PHASE_12 ? _199 : _172;
    assign _992 = ~ PHASE_12;
    assign read_enable_46 = _102 & _992;
    assign _989 = ~ _130;
    assign _990 = _129 & _989;
    assign write_enable_56 = _990 & PHASE_12;
    assign _994 = write_enable_56 | read_enable_46;
    assign address_57 = PHASE_12 ? _164 : _137;
    assign _985 = ~ PHASE_12;
    assign read_enable_47 = _102 & _985;
    assign _982 = ~ _130;
    assign _983 = _129 & _982;
    assign write_enable_57 = _983 & PHASE_12;
    assign _987 = write_enable_57 | read_enable_47;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_27
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_987), .regcea(vdd), .wea(write_enable_57), .addra(address_57), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_994), .regceb(vdd), .web(write_enable_56), .addrb(address_56), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_997[131:131]), .sbiterrb(_997[130:130]), .doutb(_997[129:66]), .dbiterra(_997[65:65]), .sbiterra(_997[64:64]), .douta(_997[63:0]) );
    assign _998 = _997[63:0];
    assign _1080 = ~ PHASE_12;
    assign _37 = _1080;
    always @(posedge _84) begin
        if (_82)
            PHASE_12 <= _980;
        else
            if (_99)
                PHASE_12 <= _37;
    end
    assign q0_3 = PHASE_12 ? _1012 : _998;
    always @(posedge _84) begin
        if (_82)
            _978 <= _977;
        else
            _978 <= _92;
    end
    assign _1069 = _978 ? _1068 : q0_3;
    dp_10
        dp_2
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1069), .d2(_1076), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1078[191:128]), .q2(_1078[127:64]), .q1(_1078[63:0]) );
    assign _1081 = _1078[63:0];
    assign data_55 = _1081;
    assign address_58 = PHASE_13 ? _164 : _68;
    assign _1145 = ~ PHASE_13;
    assign _1144 = _70[3:3];
    assign read_enable_48 = _1144 & _1145;
    always @(posedge _84) begin
        if (_82)
            _1115 <= _1114;
        else
            _1115 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1118 <= _1117;
        else
            _1118 <= _1115;
    end
    always @(posedge _84) begin
        if (_82)
            _1121 <= _1120;
        else
            _1121 <= _1118;
    end
    always @(posedge _84) begin
        if (_82)
            _1124 <= _1123;
        else
            _1124 <= _1121;
    end
    always @(posedge _84) begin
        if (_82)
            _1127 <= _1126;
        else
            _1127 <= _1124;
    end
    always @(posedge _84) begin
        if (_82)
            _1130 <= _1129;
        else
            _1130 <= _1127;
    end
    always @(posedge _84) begin
        if (_82)
            _1133 <= _1132;
        else
            _1133 <= _1130;
    end
    always @(posedge _84) begin
        if (_82)
            _1136 <= _1135;
        else
            _1136 <= _1133;
    end
    always @(posedge _84) begin
        if (_82)
            _1139 <= _1138;
        else
            _1139 <= _1136;
    end
    assign _1140 = ~ _1139;
    always @(posedge _84) begin
        if (_82)
            _1088 <= _1087;
        else
            _1088 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1091 <= _1090;
        else
            _1091 <= _1088;
    end
    always @(posedge _84) begin
        if (_82)
            _1094 <= _1093;
        else
            _1094 <= _1091;
    end
    always @(posedge _84) begin
        if (_82)
            _1097 <= _1096;
        else
            _1097 <= _1094;
    end
    always @(posedge _84) begin
        if (_82)
            _1100 <= _1099;
        else
            _1100 <= _1097;
    end
    always @(posedge _84) begin
        if (_82)
            _1103 <= _1102;
        else
            _1103 <= _1100;
    end
    always @(posedge _84) begin
        if (_82)
            _1106 <= _1105;
        else
            _1106 <= _1103;
    end
    always @(posedge _84) begin
        if (_82)
            _1109 <= _1108;
        else
            _1109 <= _1106;
    end
    always @(posedge _84) begin
        if (_82)
            _1112 <= _1111;
        else
            _1112 <= _1109;
    end
    assign _1141 = _1112 & _1140;
    assign _1142 = _129 & _1141;
    assign write_enable_58 = _1142 & PHASE_13;
    assign _1147 = write_enable_58 | read_enable_48;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_28
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1147), .regcea(vdd), .wea(write_enable_58), .addra(address_58), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_49), .regceb(vdd), .web(write_enable_49), .addrb(address_49), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1154[131:131]), .sbiterrb(_1154[130:130]), .doutb(_1154[129:66]), .dbiterra(_1154[65:65]), .sbiterra(_1154[64:64]), .douta(_1154[63:0]) );
    assign _1155 = _1154[63:0];
    assign _1085 = ~ PHASE_13;
    assign _39 = _1085;
    always @(posedge _84) begin
        if (_82)
            PHASE_13 <= _1083;
        else
            if (_72)
                PHASE_13 <= _39;
    end
    assign _1167 = PHASE_13 ? _1166 : _1155;
    assign address_59 = _1352 ? _199 : _1347;
    assign write_enable_59 = _1345 & _1352;
    assign address_60 = _1352 ? _164 : _68;
    assign _1354 = ~ _1352;
    assign read_enable_49 = _1340 & _1354;
    assign _1352 = ~ PHASE_16;
    assign write_enable_60 = _1338 & _1352;
    assign _1356 = write_enable_60 | read_enable_49;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_29
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1356), .regcea(vdd), .wea(write_enable_60), .addra(address_60), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_59), .regceb(vdd), .web(write_enable_59), .addrb(address_59), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1361[131:131]), .sbiterrb(_1361[130:130]), .doutb(_1361[129:66]), .dbiterra(_1361[65:65]), .sbiterra(_1361[64:64]), .douta(_1361[63:0]) );
    assign _1362 = _1361[63:0];
    assign address_61 = PHASE_16 ? _199 : _1347;
    assign _1345 = _129 & _1308;
    assign write_enable_61 = _1345 & PHASE_16;
    assign _1270 = _1262[129:66];
    assign _1269 = _1249[129:66];
    assign _1271 = PHASE_14 ? _1270 : _1269;
    assign _1267 = _1207[129:66];
    assign _1266 = _1193[129:66];
    assign q1_4 = PHASE_15 ? _1267 : _1266;
    assign _1272 = _1174 ? _1271 : q1_4;
    assign address_62 = _1251 ? _1245 : _1244;
    assign _1257 = ~ _1251;
    assign read_enable_50 = _102 & _1257;
    assign address_63 = _1251 ? _60 : _1227;
    assign _1253 = ~ _1251;
    assign read_enable_51 = _102 & _1253;
    assign _1251 = ~ PHASE_14;
    assign write_enable_63 = _1210 & _1251;
    assign _1255 = write_enable_63 | read_enable_51;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_30
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1255), .regcea(vdd), .wea(write_enable_63), .addra(address_63), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_50), .regceb(vdd), .web(write_enable_62), .addrb(address_62), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1262[131:131]), .sbiterrb(_1262[130:130]), .doutb(_1262[129:66]), .dbiterra(_1262[65:65]), .sbiterra(_1262[64:64]), .douta(_1262[63:0]) );
    assign _1263 = _1262[63:0];
    assign _1243 = _172[11:11];
    assign _1242 = _172[10:10];
    assign _1241 = _172[9:9];
    assign _1240 = _172[8:8];
    assign _1239 = _172[7:7];
    assign _1238 = _172[6:6];
    assign _1237 = _172[5:5];
    assign _1236 = _172[4:4];
    assign _1235 = _172[3:3];
    assign _1234 = _172[2:2];
    assign _1233 = _172[1:1];
    assign _1232 = _172[0:0];
    assign _1244 = { _1232, _1233, _1234, _1235, _1236, _1237, _1238, _1239, _1240, _1241, _1242, _1243 };
    assign address_64 = PHASE_14 ? _1245 : _1244;
    assign _1229 = ~ PHASE_14;
    assign read_enable_52 = _102 & _1229;
    assign data_61 = wr_d2;
    assign _1226 = _137[11:11];
    assign _1225 = _137[10:10];
    assign _1224 = _137[9:9];
    assign _1223 = _137[8:8];
    assign _1222 = _137[7:7];
    assign _1221 = _137[6:6];
    assign _1220 = _137[5:5];
    assign _1219 = _137[4:4];
    assign _1218 = _137[3:3];
    assign _1217 = _137[2:2];
    assign _1216 = _137[1:1];
    assign _1215 = _137[0:0];
    assign _1227 = { _1215, _1216, _1217, _1218, _1219, _1220, _1221, _1222, _1223, _1224, _1225, _1226 };
    assign address_65 = PHASE_14 ? _60 : _1227;
    assign _1212 = ~ PHASE_14;
    assign read_enable_53 = _102 & _1212;
    assign _1210 = _62[2:2];
    assign write_enable_65 = _1210 & PHASE_14;
    assign _1214 = write_enable_65 | read_enable_53;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_31
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1214), .regcea(vdd), .wea(write_enable_65), .addra(address_65), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_52), .regceb(vdd), .web(write_enable_64), .addrb(address_64), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1249[131:131]), .sbiterrb(_1249[130:130]), .doutb(_1249[129:66]), .dbiterra(_1249[65:65]), .sbiterra(_1249[64:64]), .douta(_1249[63:0]) );
    assign _1250 = _1249[63:0];
    assign _1171 = ~ PHASE_14;
    assign _43 = _1171;
    always @(posedge _84) begin
        if (_82)
            PHASE_14 <= _1169;
        else
            if (_72)
                PHASE_14 <= _43;
    end
    assign _1264 = PHASE_14 ? _1263 : _1250;
    assign address_66 = _1195 ? _199 : _172;
    assign _1202 = ~ _1195;
    assign read_enable_54 = _102 & _1202;
    assign write_enable_66 = _1186 & _1195;
    assign _1204 = write_enable_66 | read_enable_54;
    assign address_67 = _1195 ? _164 : _137;
    assign _1197 = ~ _1195;
    assign read_enable_55 = _102 & _1197;
    assign _1195 = ~ PHASE_15;
    assign write_enable_67 = _1179 & _1195;
    assign _1199 = write_enable_67 | read_enable_55;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_32
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1199), .regcea(vdd), .wea(write_enable_67), .addra(address_67), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1204), .regceb(vdd), .web(write_enable_66), .addrb(address_66), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1207[131:131]), .sbiterrb(_1207[130:130]), .doutb(_1207[129:66]), .dbiterra(_1207[65:65]), .sbiterra(_1207[64:64]), .douta(_1207[63:0]) );
    assign _1208 = _1207[63:0];
    assign _1275 = _1274[127:64];
    assign data_63 = _1275;
    assign address_68 = PHASE_15 ? _199 : _172;
    assign _1188 = ~ PHASE_15;
    assign read_enable_56 = _102 & _1188;
    assign _1185 = ~ _130;
    assign _1186 = _129 & _1185;
    assign write_enable_68 = _1186 & PHASE_15;
    assign _1190 = write_enable_68 | read_enable_56;
    assign address_69 = PHASE_15 ? _164 : _137;
    assign _1181 = ~ PHASE_15;
    assign read_enable_57 = _102 & _1181;
    assign _1178 = ~ _130;
    assign _1179 = _129 & _1178;
    assign write_enable_69 = _1179 & PHASE_15;
    assign _1183 = write_enable_69 | read_enable_57;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_33
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1183), .regcea(vdd), .wea(write_enable_69), .addra(address_69), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1190), .regceb(vdd), .web(write_enable_68), .addrb(address_68), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1193[131:131]), .sbiterrb(_1193[130:130]), .doutb(_1193[129:66]), .dbiterra(_1193[65:65]), .sbiterra(_1193[64:64]), .douta(_1193[63:0]) );
    assign _1194 = _1193[63:0];
    assign _1276 = ~ PHASE_15;
    assign _45 = _1276;
    always @(posedge _84) begin
        if (_82)
            PHASE_15 <= _1176;
        else
            if (_99)
                PHASE_15 <= _45;
    end
    assign q0_4 = PHASE_15 ? _1208 : _1194;
    always @(posedge _84) begin
        if (_82)
            _1174 <= _1173;
        else
            _1174 <= _92;
    end
    assign _1265 = _1174 ? _1264 : q0_4;
    dp_9
        dp_1
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1265), .d2(_1272), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1274[191:128]), .q2(_1274[127:64]), .q1(_1274[63:0]) );
    assign _1277 = _1274[63:0];
    assign data_67 = _1277;
    assign address_70 = PHASE_16 ? _164 : _68;
    assign _1341 = ~ PHASE_16;
    assign _1340 = _70[2:2];
    assign read_enable_58 = _1340 & _1341;
    always @(posedge _84) begin
        if (_82)
            _1311 <= _1310;
        else
            _1311 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1314 <= _1313;
        else
            _1314 <= _1311;
    end
    always @(posedge _84) begin
        if (_82)
            _1317 <= _1316;
        else
            _1317 <= _1314;
    end
    always @(posedge _84) begin
        if (_82)
            _1320 <= _1319;
        else
            _1320 <= _1317;
    end
    always @(posedge _84) begin
        if (_82)
            _1323 <= _1322;
        else
            _1323 <= _1320;
    end
    always @(posedge _84) begin
        if (_82)
            _1326 <= _1325;
        else
            _1326 <= _1323;
    end
    always @(posedge _84) begin
        if (_82)
            _1329 <= _1328;
        else
            _1329 <= _1326;
    end
    always @(posedge _84) begin
        if (_82)
            _1332 <= _1331;
        else
            _1332 <= _1329;
    end
    always @(posedge _84) begin
        if (_82)
            _1335 <= _1334;
        else
            _1335 <= _1332;
    end
    assign _1336 = ~ _1335;
    always @(posedge _84) begin
        if (_82)
            _1284 <= _1283;
        else
            _1284 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1287 <= _1286;
        else
            _1287 <= _1284;
    end
    always @(posedge _84) begin
        if (_82)
            _1290 <= _1289;
        else
            _1290 <= _1287;
    end
    always @(posedge _84) begin
        if (_82)
            _1293 <= _1292;
        else
            _1293 <= _1290;
    end
    always @(posedge _84) begin
        if (_82)
            _1296 <= _1295;
        else
            _1296 <= _1293;
    end
    always @(posedge _84) begin
        if (_82)
            _1299 <= _1298;
        else
            _1299 <= _1296;
    end
    always @(posedge _84) begin
        if (_82)
            _1302 <= _1301;
        else
            _1302 <= _1299;
    end
    always @(posedge _84) begin
        if (_82)
            _1305 <= _1304;
        else
            _1305 <= _1302;
    end
    always @(posedge _84) begin
        if (_82)
            _1308 <= _1307;
        else
            _1308 <= _1305;
    end
    assign _1337 = _1308 & _1336;
    assign _1338 = _129 & _1337;
    assign write_enable_70 = _1338 & PHASE_16;
    assign _1343 = write_enable_70 | read_enable_58;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_34
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1343), .regcea(vdd), .wea(write_enable_70), .addra(address_70), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_61), .regceb(vdd), .web(write_enable_61), .addrb(address_61), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1350[131:131]), .sbiterrb(_1350[130:130]), .doutb(_1350[129:66]), .dbiterra(_1350[65:65]), .sbiterra(_1350[64:64]), .douta(_1350[63:0]) );
    assign _1351 = _1350[63:0];
    assign _1281 = ~ PHASE_16;
    assign _47 = _1281;
    always @(posedge _84) begin
        if (_82)
            PHASE_16 <= _1279;
        else
            if (_72)
                PHASE_16 <= _47;
    end
    assign _1363 = PHASE_16 ? _1362 : _1351;
    assign address_71 = _1548 ? _199 : _1543;
    assign write_enable_71 = _1541 & _1548;
    assign address_72 = _1548 ? _164 : _68;
    assign _1550 = ~ _1548;
    assign read_enable_59 = _1536 & _1550;
    assign _1548 = ~ PHASE_19;
    assign write_enable_72 = _1534 & _1548;
    assign _1552 = write_enable_72 | read_enable_59;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_35
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1552), .regcea(vdd), .wea(write_enable_72), .addra(address_72), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_71), .regceb(vdd), .web(write_enable_71), .addrb(address_71), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1557[131:131]), .sbiterrb(_1557[130:130]), .doutb(_1557[129:66]), .dbiterra(_1557[65:65]), .sbiterra(_1557[64:64]), .douta(_1557[63:0]) );
    assign _1558 = _1557[63:0];
    assign address_73 = PHASE_19 ? _199 : _1543;
    assign _1541 = _129 & _1504;
    assign write_enable_73 = _1541 & PHASE_19;
    assign _1466 = _1458[129:66];
    assign _1465 = _1445[129:66];
    assign _1467 = PHASE_17 ? _1466 : _1465;
    assign _1463 = _1403[129:66];
    assign _1462 = _1389[129:66];
    assign q1_5 = PHASE_18 ? _1463 : _1462;
    assign _1468 = _1370 ? _1467 : q1_5;
    assign address_74 = _1447 ? _1441 : _1440;
    assign _1453 = ~ _1447;
    assign read_enable_60 = _102 & _1453;
    assign address_75 = _1447 ? _60 : _1423;
    assign _1449 = ~ _1447;
    assign read_enable_61 = _102 & _1449;
    assign _1447 = ~ PHASE_17;
    assign write_enable_75 = _1406 & _1447;
    assign _1451 = write_enable_75 | read_enable_61;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_36
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1451), .regcea(vdd), .wea(write_enable_75), .addra(address_75), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_60), .regceb(vdd), .web(write_enable_74), .addrb(address_74), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1458[131:131]), .sbiterrb(_1458[130:130]), .doutb(_1458[129:66]), .dbiterra(_1458[65:65]), .sbiterra(_1458[64:64]), .douta(_1458[63:0]) );
    assign _1459 = _1458[63:0];
    assign _1439 = _172[11:11];
    assign _1438 = _172[10:10];
    assign _1437 = _172[9:9];
    assign _1436 = _172[8:8];
    assign _1435 = _172[7:7];
    assign _1434 = _172[6:6];
    assign _1433 = _172[5:5];
    assign _1432 = _172[4:4];
    assign _1431 = _172[3:3];
    assign _1430 = _172[2:2];
    assign _1429 = _172[1:1];
    assign _1428 = _172[0:0];
    assign _1440 = { _1428, _1429, _1430, _1431, _1432, _1433, _1434, _1435, _1436, _1437, _1438, _1439 };
    assign address_76 = PHASE_17 ? _1441 : _1440;
    assign _1425 = ~ PHASE_17;
    assign read_enable_62 = _102 & _1425;
    assign data_73 = wr_d1;
    assign _1422 = _137[11:11];
    assign _1421 = _137[10:10];
    assign _1420 = _137[9:9];
    assign _1419 = _137[8:8];
    assign _1418 = _137[7:7];
    assign _1417 = _137[6:6];
    assign _1416 = _137[5:5];
    assign _1415 = _137[4:4];
    assign _1414 = _137[3:3];
    assign _1413 = _137[2:2];
    assign _1412 = _137[1:1];
    assign _1411 = _137[0:0];
    assign _1423 = { _1411, _1412, _1413, _1414, _1415, _1416, _1417, _1418, _1419, _1420, _1421, _1422 };
    assign address_77 = PHASE_17 ? _60 : _1423;
    assign _1408 = ~ PHASE_17;
    assign read_enable_63 = _102 & _1408;
    assign _1406 = _62[1:1];
    assign write_enable_77 = _1406 & PHASE_17;
    assign _1410 = write_enable_77 | read_enable_63;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_37
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1410), .regcea(vdd), .wea(write_enable_77), .addra(address_77), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_62), .regceb(vdd), .web(write_enable_76), .addrb(address_76), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1445[131:131]), .sbiterrb(_1445[130:130]), .doutb(_1445[129:66]), .dbiterra(_1445[65:65]), .sbiterra(_1445[64:64]), .douta(_1445[63:0]) );
    assign _1446 = _1445[63:0];
    assign _1367 = ~ PHASE_17;
    assign _51 = _1367;
    always @(posedge _84) begin
        if (_82)
            PHASE_17 <= _1365;
        else
            if (_72)
                PHASE_17 <= _51;
    end
    assign _1460 = PHASE_17 ? _1459 : _1446;
    assign address_78 = _1391 ? _199 : _172;
    assign _1398 = ~ _1391;
    assign read_enable_64 = _102 & _1398;
    assign write_enable_78 = _1382 & _1391;
    assign _1400 = write_enable_78 | read_enable_64;
    assign address_79 = _1391 ? _164 : _137;
    assign _1393 = ~ _1391;
    assign read_enable_65 = _102 & _1393;
    assign _1391 = ~ PHASE_18;
    assign write_enable_79 = _1375 & _1391;
    assign _1395 = write_enable_79 | read_enable_65;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_38
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1395), .regcea(vdd), .wea(write_enable_79), .addra(address_79), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1400), .regceb(vdd), .web(write_enable_78), .addrb(address_78), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1403[131:131]), .sbiterrb(_1403[130:130]), .doutb(_1403[129:66]), .dbiterra(_1403[65:65]), .sbiterra(_1403[64:64]), .douta(_1403[63:0]) );
    assign _1404 = _1403[63:0];
    assign _1471 = _1470[127:64];
    assign data_75 = _1471;
    assign address_80 = PHASE_18 ? _199 : _172;
    assign _1384 = ~ PHASE_18;
    assign read_enable_66 = _102 & _1384;
    assign _1381 = ~ _130;
    assign _1382 = _129 & _1381;
    assign write_enable_80 = _1382 & PHASE_18;
    assign _1386 = write_enable_80 | read_enable_66;
    assign address_81 = PHASE_18 ? _164 : _137;
    assign _1377 = ~ PHASE_18;
    assign read_enable_67 = _102 & _1377;
    assign _1374 = ~ _130;
    assign _1375 = _129 & _1374;
    assign write_enable_81 = _1375 & PHASE_18;
    assign _1379 = write_enable_81 | read_enable_67;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_39
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1379), .regcea(vdd), .wea(write_enable_81), .addra(address_81), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1386), .regceb(vdd), .web(write_enable_80), .addrb(address_80), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1389[131:131]), .sbiterrb(_1389[130:130]), .doutb(_1389[129:66]), .dbiterra(_1389[65:65]), .sbiterra(_1389[64:64]), .douta(_1389[63:0]) );
    assign _1390 = _1389[63:0];
    assign _1472 = ~ PHASE_18;
    assign _53 = _1472;
    always @(posedge _84) begin
        if (_82)
            PHASE_18 <= _1372;
        else
            if (_99)
                PHASE_18 <= _53;
    end
    assign q0_5 = PHASE_18 ? _1404 : _1390;
    always @(posedge _84) begin
        if (_82)
            _1370 <= _1369;
        else
            _1370 <= _92;
    end
    assign _1461 = _1370 ? _1460 : q0_5;
    dp_8
        dp_0
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1461), .d2(_1468), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1470[191:128]), .q2(_1470[127:64]), .q1(_1470[63:0]) );
    assign _1473 = _1470[63:0];
    assign data_79 = _1473;
    assign address_82 = PHASE_19 ? _164 : _68;
    assign _1537 = ~ PHASE_19;
    assign _1536 = _70[1:1];
    assign read_enable_68 = _1536 & _1537;
    always @(posedge _84) begin
        if (_82)
            _1507 <= _1506;
        else
            _1507 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1510 <= _1509;
        else
            _1510 <= _1507;
    end
    always @(posedge _84) begin
        if (_82)
            _1513 <= _1512;
        else
            _1513 <= _1510;
    end
    always @(posedge _84) begin
        if (_82)
            _1516 <= _1515;
        else
            _1516 <= _1513;
    end
    always @(posedge _84) begin
        if (_82)
            _1519 <= _1518;
        else
            _1519 <= _1516;
    end
    always @(posedge _84) begin
        if (_82)
            _1522 <= _1521;
        else
            _1522 <= _1519;
    end
    always @(posedge _84) begin
        if (_82)
            _1525 <= _1524;
        else
            _1525 <= _1522;
    end
    always @(posedge _84) begin
        if (_82)
            _1528 <= _1527;
        else
            _1528 <= _1525;
    end
    always @(posedge _84) begin
        if (_82)
            _1531 <= _1530;
        else
            _1531 <= _1528;
    end
    assign _1532 = ~ _1531;
    always @(posedge _84) begin
        if (_82)
            _1480 <= _1479;
        else
            _1480 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1483 <= _1482;
        else
            _1483 <= _1480;
    end
    always @(posedge _84) begin
        if (_82)
            _1486 <= _1485;
        else
            _1486 <= _1483;
    end
    always @(posedge _84) begin
        if (_82)
            _1489 <= _1488;
        else
            _1489 <= _1486;
    end
    always @(posedge _84) begin
        if (_82)
            _1492 <= _1491;
        else
            _1492 <= _1489;
    end
    always @(posedge _84) begin
        if (_82)
            _1495 <= _1494;
        else
            _1495 <= _1492;
    end
    always @(posedge _84) begin
        if (_82)
            _1498 <= _1497;
        else
            _1498 <= _1495;
    end
    always @(posedge _84) begin
        if (_82)
            _1501 <= _1500;
        else
            _1501 <= _1498;
    end
    always @(posedge _84) begin
        if (_82)
            _1504 <= _1503;
        else
            _1504 <= _1501;
    end
    assign _1533 = _1504 & _1532;
    assign _1534 = _129 & _1533;
    assign write_enable_82 = _1534 & PHASE_19;
    assign _1539 = write_enable_82 | read_enable_68;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_40
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1539), .regcea(vdd), .wea(write_enable_82), .addra(address_82), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_73), .regceb(vdd), .web(write_enable_73), .addrb(address_73), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1546[131:131]), .sbiterrb(_1546[130:130]), .doutb(_1546[129:66]), .dbiterra(_1546[65:65]), .sbiterra(_1546[64:64]), .douta(_1546[63:0]) );
    assign _1547 = _1546[63:0];
    assign _1477 = ~ PHASE_19;
    assign _55 = _1477;
    always @(posedge _84) begin
        if (_82)
            PHASE_19 <= _1475;
        else
            if (_72)
                PHASE_19 <= _55;
    end
    assign _1559 = PHASE_19 ? _1558 : _1547;
    assign address_83 = _1744 ? _199 : _1739;
    assign write_enable_83 = _1737 & _1744;
    assign address_84 = _1744 ? _164 : _68;
    assign _1746 = ~ _1744;
    assign read_enable_69 = _1732 & _1746;
    assign _1744 = ~ PHASE_22;
    assign write_enable_84 = _1730 & _1744;
    assign _1748 = write_enable_84 | read_enable_69;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_41
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1748), .regcea(vdd), .wea(write_enable_84), .addra(address_84), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_83), .regceb(vdd), .web(write_enable_83), .addrb(address_83), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1753[131:131]), .sbiterrb(_1753[130:130]), .doutb(_1753[129:66]), .dbiterra(_1753[65:65]), .sbiterra(_1753[64:64]), .douta(_1753[63:0]) );
    assign _1754 = _1753[63:0];
    assign address_85 = PHASE_22 ? _199 : _1739;
    assign _1737 = _129 & _1700;
    assign write_enable_85 = _1737 & PHASE_22;
    assign _292 = _91[521:518];
    assign _291 = _91[517:517];
    assign _289 = _91[513:513];
    assign _288 = _91[512:449];
    assign _287 = _91[448:385];
    assign _286 = _91[384:321];
    assign _285 = _91[320:257];
    assign _284 = _91[256:193];
    assign _283 = _91[192:129];
    assign _282 = _91[128:65];
    assign _1662 = _1654[129:66];
    assign _1661 = _1641[129:66];
    assign _1663 = PHASE_20 ? _1662 : _1661;
    assign _1659 = _1599[129:66];
    assign _1658 = _1585[129:66];
    assign q1_6 = PHASE_21 ? _1659 : _1658;
    assign _1664 = _1566 ? _1663 : q1_6;
    assign address_86 = _1643 ? _1637 : _1636;
    assign _1649 = ~ _1643;
    assign read_enable_70 = _102 & _1649;
    assign address_87 = _1643 ? _60 : _1619;
    assign _1645 = ~ _1643;
    assign read_enable_71 = _102 & _1645;
    assign _1643 = ~ PHASE_20;
    assign write_enable_87 = _1602 & _1643;
    assign _1647 = write_enable_87 | read_enable_71;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_42
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1647), .regcea(vdd), .wea(write_enable_87), .addra(address_87), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_70), .regceb(vdd), .web(write_enable_86), .addrb(address_86), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1654[131:131]), .sbiterrb(_1654[130:130]), .doutb(_1654[129:66]), .dbiterra(_1654[65:65]), .sbiterra(_1654[64:64]), .douta(_1654[63:0]) );
    assign _1655 = _1654[63:0];
    assign _1635 = _172[11:11];
    assign _1634 = _172[10:10];
    assign _1633 = _172[9:9];
    assign _1632 = _172[8:8];
    assign _1631 = _172[7:7];
    assign _1630 = _172[6:6];
    assign _1629 = _172[5:5];
    assign _1628 = _172[4:4];
    assign _1627 = _172[3:3];
    assign _1626 = _172[2:2];
    assign _1625 = _172[1:1];
    assign _1624 = _172[0:0];
    assign _1636 = { _1624, _1625, _1626, _1627, _1628, _1629, _1630, _1631, _1632, _1633, _1634, _1635 };
    assign address_88 = PHASE_20 ? _1637 : _1636;
    assign _1621 = ~ PHASE_20;
    assign read_enable_72 = _102 & _1621;
    assign data_85 = wr_d0;
    assign _60 = wr_addr;
    assign _1618 = _137[11:11];
    assign _1617 = _137[10:10];
    assign _1616 = _137[9:9];
    assign _1615 = _137[8:8];
    assign _1614 = _137[7:7];
    assign _1613 = _137[6:6];
    assign _1612 = _137[5:5];
    assign _1611 = _137[4:4];
    assign _1610 = _137[3:3];
    assign _1609 = _137[2:2];
    assign _1608 = _137[1:1];
    assign _1607 = _137[0:0];
    assign _1619 = { _1607, _1608, _1609, _1610, _1611, _1612, _1613, _1614, _1615, _1616, _1617, _1618 };
    assign address_89 = PHASE_20 ? _60 : _1619;
    assign _1604 = ~ PHASE_20;
    assign read_enable_73 = _102 & _1604;
    assign _62 = wr_en;
    assign _1602 = _62[0:0];
    assign write_enable_89 = _1602 & PHASE_20;
    assign _1606 = write_enable_89 | read_enable_73;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_43
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1606), .regcea(vdd), .wea(write_enable_89), .addra(address_89), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_72), .regceb(vdd), .web(write_enable_88), .addrb(address_88), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1641[131:131]), .sbiterrb(_1641[130:130]), .doutb(_1641[129:66]), .dbiterra(_1641[65:65]), .sbiterra(_1641[64:64]), .douta(_1641[63:0]) );
    assign _1642 = _1641[63:0];
    assign _1563 = ~ PHASE_20;
    assign _63 = _1563;
    always @(posedge _84) begin
        if (_82)
            PHASE_20 <= _1561;
        else
            if (_72)
                PHASE_20 <= _63;
    end
    assign _1656 = PHASE_20 ? _1655 : _1642;
    assign address_90 = _1587 ? _199 : _172;
    assign _1594 = ~ _1587;
    assign read_enable_74 = _102 & _1594;
    assign write_enable_90 = _1578 & _1587;
    assign _1596 = write_enable_90 | read_enable_74;
    assign address_91 = _1587 ? _164 : _137;
    assign _1589 = ~ _1587;
    assign read_enable_75 = _102 & _1589;
    assign _1587 = ~ PHASE_21;
    assign write_enable_91 = _1571 & _1587;
    assign _1591 = write_enable_91 | read_enable_75;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_44
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1591), .regcea(vdd), .wea(write_enable_91), .addra(address_91), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1596), .regceb(vdd), .web(write_enable_90), .addrb(address_90), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1599[131:131]), .sbiterrb(_1599[130:130]), .doutb(_1599[129:66]), .dbiterra(_1599[65:65]), .sbiterra(_1599[64:64]), .douta(_1599[63:0]) );
    assign _1600 = _1599[63:0];
    assign _1667 = _1666[127:64];
    assign data_87 = _1667;
    always @(posedge _84) begin
        if (_82)
            _175 <= _174;
        else
            _175 <= _172;
    end
    always @(posedge _84) begin
        if (_82)
            _178 <= _177;
        else
            _178 <= _175;
    end
    always @(posedge _84) begin
        if (_82)
            _181 <= _180;
        else
            _181 <= _178;
    end
    always @(posedge _84) begin
        if (_82)
            _184 <= _183;
        else
            _184 <= _181;
    end
    always @(posedge _84) begin
        if (_82)
            _187 <= _186;
        else
            _187 <= _184;
    end
    always @(posedge _84) begin
        if (_82)
            _190 <= _189;
        else
            _190 <= _187;
    end
    always @(posedge _84) begin
        if (_82)
            _193 <= _192;
        else
            _193 <= _190;
    end
    always @(posedge _84) begin
        if (_82)
            _196 <= _195;
        else
            _196 <= _193;
    end
    always @(posedge _84) begin
        if (_82)
            _199 <= _198;
        else
            _199 <= _196;
    end
    assign _172 = _91[64:53];
    assign address_92 = PHASE_21 ? _199 : _172;
    assign _1580 = ~ PHASE_21;
    assign read_enable_76 = _102 & _1580;
    assign _1577 = ~ _130;
    assign _1578 = _129 & _1577;
    assign write_enable_92 = _1578 & PHASE_21;
    assign _1582 = write_enable_92 | read_enable_76;
    assign address_93 = PHASE_21 ? _164 : _137;
    assign _1573 = ~ PHASE_21;
    assign read_enable_77 = _102 & _1573;
    assign _1570 = ~ _130;
    assign _1571 = _129 & _1570;
    assign write_enable_93 = _1571 & PHASE_21;
    assign _1575 = write_enable_93 | read_enable_77;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_45
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1575), .regcea(vdd), .wea(write_enable_93), .addra(address_93), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1582), .regceb(vdd), .web(write_enable_92), .addrb(address_92), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1585[131:131]), .sbiterrb(_1585[130:130]), .doutb(_1585[129:66]), .dbiterra(_1585[65:65]), .sbiterra(_1585[64:64]), .douta(_1585[63:0]) );
    assign _1586 = _1585[63:0];
    assign _99 = _91[523:523];
    assign _1668 = ~ PHASE_21;
    assign _65 = _1668;
    always @(posedge _84) begin
        if (_82)
            PHASE_21 <= _1568;
        else
            if (_99)
                PHASE_21 <= _65;
    end
    assign q0_6 = PHASE_21 ? _1600 : _1586;
    assign _92 = _91[514:514];
    always @(posedge _84) begin
        if (_82)
            _1566 <= _1565;
        else
            _1566 <= _92;
    end
    assign _1657 = _1566 ? _1656 : q0_6;
    dp_7
        dp
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1657), .d2(_1664), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1666[191:128]), .q2(_1666[127:64]), .q1(_1666[63:0]) );
    assign _1669 = _1666[63:0];
    assign data_91 = _1669;
    assign _137 = _91[52:41];
    always @(posedge _84) begin
        if (_82)
            _140 <= _139;
        else
            _140 <= _137;
    end
    always @(posedge _84) begin
        if (_82)
            _143 <= _142;
        else
            _143 <= _140;
    end
    always @(posedge _84) begin
        if (_82)
            _146 <= _145;
        else
            _146 <= _143;
    end
    always @(posedge _84) begin
        if (_82)
            _149 <= _148;
        else
            _149 <= _146;
    end
    always @(posedge _84) begin
        if (_82)
            _152 <= _151;
        else
            _152 <= _149;
    end
    always @(posedge _84) begin
        if (_82)
            _155 <= _154;
        else
            _155 <= _152;
    end
    always @(posedge _84) begin
        if (_82)
            _158 <= _157;
        else
            _158 <= _155;
    end
    always @(posedge _84) begin
        if (_82)
            _161 <= _160;
        else
            _161 <= _158;
    end
    always @(posedge _84) begin
        if (_82)
            _164 <= _163;
        else
            _164 <= _161;
    end
    assign _68 = rd_addr;
    assign address_94 = PHASE_22 ? _164 : _68;
    assign _1733 = ~ PHASE_22;
    assign _70 = rd_en;
    assign _1732 = _70[0:0];
    assign read_enable_78 = _1732 & _1733;
    assign _290 = _91[516:516];
    always @(posedge _84) begin
        if (_82)
            _1703 <= _1702;
        else
            _1703 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1706 <= _1705;
        else
            _1706 <= _1703;
    end
    always @(posedge _84) begin
        if (_82)
            _1709 <= _1708;
        else
            _1709 <= _1706;
    end
    always @(posedge _84) begin
        if (_82)
            _1712 <= _1711;
        else
            _1712 <= _1709;
    end
    always @(posedge _84) begin
        if (_82)
            _1715 <= _1714;
        else
            _1715 <= _1712;
    end
    always @(posedge _84) begin
        if (_82)
            _1718 <= _1717;
        else
            _1718 <= _1715;
    end
    always @(posedge _84) begin
        if (_82)
            _1721 <= _1720;
        else
            _1721 <= _1718;
    end
    always @(posedge _84) begin
        if (_82)
            _1724 <= _1723;
        else
            _1724 <= _1721;
    end
    always @(posedge _84) begin
        if (_82)
            _1727 <= _1726;
        else
            _1727 <= _1724;
    end
    assign _1728 = ~ _1727;
    assign _130 = _91[515:515];
    always @(posedge _84) begin
        if (_82)
            _1676 <= _1675;
        else
            _1676 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1679 <= _1678;
        else
            _1679 <= _1676;
    end
    always @(posedge _84) begin
        if (_82)
            _1682 <= _1681;
        else
            _1682 <= _1679;
    end
    always @(posedge _84) begin
        if (_82)
            _1685 <= _1684;
        else
            _1685 <= _1682;
    end
    always @(posedge _84) begin
        if (_82)
            _1688 <= _1687;
        else
            _1688 <= _1685;
    end
    always @(posedge _84) begin
        if (_82)
            _1691 <= _1690;
        else
            _1691 <= _1688;
    end
    always @(posedge _84) begin
        if (_82)
            _1694 <= _1693;
        else
            _1694 <= _1691;
    end
    always @(posedge _84) begin
        if (_82)
            _1697 <= _1696;
        else
            _1697 <= _1694;
    end
    always @(posedge _84) begin
        if (_82)
            _1700 <= _1699;
        else
            _1700 <= _1697;
    end
    assign _1729 = _1700 & _1728;
    assign _102 = _91[522:522];
    always @(posedge _84) begin
        if (_82)
            _105 <= _104;
        else
            _105 <= _102;
    end
    always @(posedge _84) begin
        if (_82)
            _108 <= _107;
        else
            _108 <= _105;
    end
    always @(posedge _84) begin
        if (_82)
            _111 <= _110;
        else
            _111 <= _108;
    end
    always @(posedge _84) begin
        if (_82)
            _114 <= _113;
        else
            _114 <= _111;
    end
    always @(posedge _84) begin
        if (_82)
            _117 <= _116;
        else
            _117 <= _114;
    end
    always @(posedge _84) begin
        if (_82)
            _120 <= _119;
        else
            _120 <= _117;
    end
    always @(posedge _84) begin
        if (_82)
            _123 <= _122;
        else
            _123 <= _120;
    end
    always @(posedge _84) begin
        if (_82)
            _126 <= _125;
        else
            _126 <= _123;
    end
    always @(posedge _84) begin
        if (_82)
            _129 <= _128;
        else
            _129 <= _126;
    end
    assign _1730 = _129 & _1729;
    assign write_enable_94 = _1730 & PHASE_22;
    assign _1735 = write_enable_94 | read_enable_78;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_46
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1735), .regcea(vdd), .wea(write_enable_94), .addra(address_94), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_85), .regceb(vdd), .web(write_enable_85), .addrb(address_85), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1742[131:131]), .sbiterrb(_1742[130:130]), .doutb(_1742[129:66]), .dbiterra(_1742[65:65]), .sbiterra(_1742[64:64]), .douta(_1742[63:0]) );
    assign _1743 = _1742[63:0];
    assign _72 = flip;
    assign _1673 = ~ PHASE_22;
    assign _73 = _1673;
    always @(posedge _84) begin
        if (_82)
            PHASE_22 <= _1671;
        else
            if (_72)
                PHASE_22 <= _73;
    end
    assign _1755 = PHASE_22 ? _1754 : _1743;
    assign _76 = first_4step_pass;
    assign _78 = first_iter;
    assign _80 = start;
    assign _82 = clear;
    assign _84 = clock;
    ctrl
        ctrl
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .first_4step_pass(_76), .flip(_91[523:523]), .read_write_enable(_91[522:522]), .index(_91[521:518]), .valid(_91[517:517]), .twiddle_stage(_91[516:516]), .last_stage(_91[515:515]), .first_stage(_91[514:514]), .start_twiddles(_91[513:513]), .omegas6(_91[512:449]), .omegas5(_91[448:385]), .omegas4(_91[384:321]), .omegas3(_91[320:257]), .omegas2(_91[256:193]), .omegas1(_91[192:129]), .omegas0(_91[128:65]), .addr2(_91[64:53]), .addr1(_91[52:41]), .m(_91[40:29]), .k(_91[28:17]), .j(_91[16:5]), .i(_91[4:1]), .done_(_91[0:0]) );
    assign _1756 = _91[0:0];

    /* aliases */
    assign data_0 = data;
    assign data_2 = data_1;
    assign data_4 = data_3;
    assign data_5 = data_3;
    assign data_6 = data_3;
    assign data_8 = data_7;
    assign data_9 = data_7;
    assign data_10 = data_7;
    assign data_12 = data_11;
    assign data_14 = data_13;
    assign data_16 = data_15;
    assign data_17 = data_15;
    assign data_18 = data_15;
    assign data_20 = data_19;
    assign data_21 = data_19;
    assign data_22 = data_19;
    assign data_24 = data_23;
    assign data_26 = data_25;
    assign data_28 = data_27;
    assign data_29 = data_27;
    assign data_30 = data_27;
    assign data_32 = data_31;
    assign data_33 = data_31;
    assign data_34 = data_31;
    assign data_36 = data_35;
    assign data_38 = data_37;
    assign data_40 = data_39;
    assign data_41 = data_39;
    assign data_42 = data_39;
    assign data_44 = data_43;
    assign data_45 = data_43;
    assign data_46 = data_43;
    assign data_48 = data_47;
    assign data_50 = data_49;
    assign data_52 = data_51;
    assign data_53 = data_51;
    assign data_54 = data_51;
    assign data_56 = data_55;
    assign data_57 = data_55;
    assign data_58 = data_55;
    assign data_60 = data_59;
    assign data_62 = data_61;
    assign data_64 = data_63;
    assign data_65 = data_63;
    assign data_66 = data_63;
    assign data_68 = data_67;
    assign data_69 = data_67;
    assign data_70 = data_67;
    assign data_72 = data_71;
    assign data_74 = data_73;
    assign data_76 = data_75;
    assign data_77 = data_75;
    assign data_78 = data_75;
    assign data_80 = data_79;
    assign data_81 = data_79;
    assign data_82 = data_79;
    assign data_84 = data_83;
    assign data_86 = data_85;
    assign data_88 = data_87;
    assign data_89 = data_87;
    assign data_90 = data_87;
    assign data_92 = data_91;
    assign data_93 = data_91;
    assign data_94 = data_91;

    /* output assignments */
    assign done_ = _1756;
    assign rd_q0 = _1755;
    assign rd_q1 = _1559;
    assign rd_q2 = _1363;
    assign rd_q3 = _1167;
    assign rd_q4 = _971;
    assign rd_q5 = _775;
    assign rd_q6 = _579;
    assign rd_q7 = _383;

endmodule
module dp_15 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0001011010011001110010100011110011001100000000011000111101010101;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0110100110010111111010001101100011001001101111010100100000100101;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0010000100011110110101100011101101010010011110100001110000110111;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0000101011001010001100100100101101011011001100100000011011011100;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1111101111010100000111000110101110001100101010100011001100000010;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0011000010111010001011101100110101011110100100111110011101101101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_16 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0001111011110111101001011100000111101100100110110000000100100111;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0111111010110111000101110011011011100010101100111010000100000110;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1111000000111100000010001100010110100010100001001001001111111101;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1001110001100101101001000011100011101100100110101001011111111000;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0110000010001000010110101101110010000100111001101000101001111110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0110101111000000010111100100011101010101010001100110100011000010;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0000001100000000101001011101111000101110111111100011110111000001;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_17 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1110000101110100011000000100000100110100000010000010100100010011;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0001001000111000010111110001101011011001000001111111010110000000;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0100000110110111010100110011011100010101000101100000000101100101;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0000000110011111011011110111001101111001110110010011010011110001;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0000000010100111001011000000010010100111011101011111110001111000;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0110110010110000111011001100000000010111101011101101100010111100;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1111011001111000001001110011001110101011000101110000100110010000;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_18 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0001000110111000101011101001011001111100100001000010010100110010;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1100100010110010000000011011001100000010111000101000000110010110;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1011010100001110001010100010011100101100010010111001100001111111;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0100100010101101111000110100110001111001100110001001111000111111;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1000101010000001010100111101100011011111111101101100100000001101;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1011001111101011010100101110010011000101101010010001011100000111;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0000111010000001010111111000011100011101110010011110011101011100;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_19 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1000000000010101010101101101000101010110000010111110001110111000;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0101001110010000111001101101001110111101111110001100111010111111;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0001011111010001110111110010100111110100110100010110100100111010;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0010000100011110110101100011101101010010011110100001110000110111;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0101100000001101011100101110110101101100101000101100101011001111;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1100111100000101001110011010010101001111101000110101101001010101;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1100101111011100100111001010001111010111100111010001110111111011;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_20 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0101000011001111001101110000000110110101011011100101101000110110;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1110000101110100011000000100000100110100000010000010100100010011;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0101110100110000000100110101011101000010111111000111010000001011;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0110001110111000011110101101110010111010001011110110000001100110;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0000010100100101000010101011110010110110000000011111001101101000;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0010101001001000011111010001011101101011111100000111111100100010;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0111010000100110001111001000111100111011110010111011011011111001;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_21 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1010101010110111010011110011111010111101100110101001001011011011;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0100011111101001000011110000001000111010101011110101010100100101;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1001010100101001000110000101000110101101100000000110001101010110;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1100101000011000110011110101000000110000010010010011001010001001;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0110100101101111110010001001101110011101101001011110000011100001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1101101000101011101011101011110001010010100001010000110110101000;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1100100111010010110100011100111101011011010100100100011110000101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_22 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0100011011100001001000010000000001111110000000001111000110100011;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0001011011010010100001100000100011010110001111011101101100101001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1011001100010011101001011101010111010001000111001110100000000110;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0001001001101101010000000010001001100101110100000011001111101011;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1110011100101010111000001110100001011010010101001011001011111110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1010110100011111111111000101110001001001010010010001100001101110;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1100011000010110000110000001000110110010011000110111100111111101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module parallel_cores_1 (
    wr_d7,
    wr_d6,
    wr_d5,
    wr_d4,
    wr_d3,
    wr_d2,
    wr_d1,
    wr_d0,
    wr_addr,
    wr_en,
    rd_addr,
    rd_en,
    flip,
    first_4step_pass,
    first_iter,
    start,
    clear,
    clock,
    done_,
    rd_q0,
    rd_q1,
    rd_q2,
    rd_q3,
    rd_q4,
    rd_q5,
    rd_q6,
    rd_q7
);

    input [63:0] wr_d7;
    input [63:0] wr_d6;
    input [63:0] wr_d5;
    input [63:0] wr_d4;
    input [63:0] wr_d3;
    input [63:0] wr_d2;
    input [63:0] wr_d1;
    input [63:0] wr_d0;
    input [11:0] wr_addr;
    input [7:0] wr_en;
    input [11:0] rd_addr;
    input [7:0] rd_en;
    input flip;
    input first_4step_pass;
    input first_iter;
    input start;
    input clear;
    input clock;
    output done_;
    output [63:0] rd_q0;
    output [63:0] rd_q1;
    output [63:0] rd_q2;
    output [63:0] rd_q3;
    output [63:0] rd_q4;
    output [63:0] rd_q5;
    output [63:0] rd_q6;
    output [63:0] rd_q7;

    /* signal declarations */
    wire [11:0] address;
    wire write_enable;
    wire [11:0] address_0;
    wire _374;
    wire read_enable;
    wire _372;
    wire write_enable_0;
    wire _376;
    wire [131:0] _381;
    wire [63:0] _382;
    wire [11:0] _367 = 12'b000000000000;
    wire [11:0] address_1;
    wire _365;
    wire write_enable_1;
    wire [63:0] _279;
    wire [63:0] _278;
    wire [63:0] _280;
    wire [63:0] _276;
    wire [63:0] _275;
    wire [63:0] q1;
    wire [63:0] _281;
    wire [11:0] address_2;
    wire write_enable_2 = 1'b0;
    wire _266;
    wire read_enable_0;
    wire [11:0] address_3;
    wire _262;
    wire read_enable_1;
    wire _260;
    wire write_enable_3;
    wire _264;
    wire [131:0] _271;
    wire [63:0] _272;
    wire [63:0] data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_0;
    wire [11:0] _254 = 12'b000000000000;
    wire _252;
    wire _251;
    wire _250;
    wire _249;
    wire _248;
    wire _247;
    wire _246;
    wire _245;
    wire _244;
    wire _243;
    wire _242;
    wire _241;
    wire [11:0] _253;
    wire [11:0] address_4;
    wire write_enable_4 = 1'b0;
    wire _238;
    wire read_enable_2;
    wire [63:0] data_1;
    wire [63:0] data_2;
    wire _235;
    wire _234;
    wire _233;
    wire _232;
    wire _231;
    wire _230;
    wire _229;
    wire _228;
    wire _227;
    wire _226;
    wire _225;
    wire _224;
    wire [11:0] _236;
    wire [11:0] address_5;
    wire _221;
    wire read_enable_3;
    wire _219;
    wire write_enable_5;
    wire _223;
    wire [131:0] _258;
    wire [63:0] _259;
    wire _87 = 1'b0;
    wire _86 = 1'b0;
    wire _89;
    wire _3;
    reg PHASE;
    wire [63:0] _273;
    wire [11:0] address_6;
    wire _211;
    wire read_enable_4;
    wire write_enable_6;
    wire _213;
    wire [11:0] address_7;
    wire _206;
    wire read_enable_5;
    wire _204;
    wire write_enable_7;
    wire _208;
    wire [131:0] _216;
    wire [63:0] _217;
    wire [63:0] _295;
    wire [63:0] data_3;
    wire [63:0] data_4;
    wire [63:0] data_5;
    wire [63:0] data_6;
    wire [11:0] address_8;
    wire _169;
    wire read_enable_6;
    wire _166;
    wire _167;
    wire write_enable_8;
    wire _171;
    wire [11:0] address_9;
    wire _134;
    wire read_enable_7;
    wire _131;
    wire _132;
    wire write_enable_9;
    wire _136;
    wire [131:0] _202;
    wire [63:0] _203;
    wire _98 = 1'b0;
    wire _97 = 1'b0;
    wire _296;
    wire _5;
    reg PHASE_0;
    wire [63:0] q0;
    wire _94 = 1'b0;
    wire _93 = 1'b0;
    reg _96;
    wire [63:0] _274;
    wire [191:0] _294;
    wire [63:0] _297;
    wire [63:0] data_7;
    wire [63:0] data_8;
    wire [63:0] data_9;
    wire [63:0] data_10;
    wire [11:0] address_10;
    wire _361;
    wire _360;
    wire read_enable_8;
    wire _354 = 1'b0;
    wire _353 = 1'b0;
    wire _351 = 1'b0;
    wire _350 = 1'b0;
    wire _348 = 1'b0;
    wire _347 = 1'b0;
    wire _345 = 1'b0;
    wire _344 = 1'b0;
    wire _342 = 1'b0;
    wire _341 = 1'b0;
    wire _339 = 1'b0;
    wire _338 = 1'b0;
    wire _336 = 1'b0;
    wire _335 = 1'b0;
    wire _333 = 1'b0;
    wire _332 = 1'b0;
    wire _330 = 1'b0;
    wire _329 = 1'b0;
    reg _331;
    reg _334;
    reg _337;
    reg _340;
    reg _343;
    reg _346;
    reg _349;
    reg _352;
    reg _355;
    wire _356;
    wire _327 = 1'b0;
    wire _326 = 1'b0;
    wire _324 = 1'b0;
    wire _323 = 1'b0;
    wire _321 = 1'b0;
    wire _320 = 1'b0;
    wire _318 = 1'b0;
    wire _317 = 1'b0;
    wire _315 = 1'b0;
    wire _314 = 1'b0;
    wire _312 = 1'b0;
    wire _311 = 1'b0;
    wire _309 = 1'b0;
    wire _308 = 1'b0;
    wire _306 = 1'b0;
    wire _305 = 1'b0;
    wire _303 = 1'b0;
    wire _302 = 1'b0;
    reg _304;
    reg _307;
    reg _310;
    reg _313;
    reg _316;
    reg _319;
    reg _322;
    reg _325;
    reg _328;
    wire _357;
    wire _358;
    wire write_enable_10;
    wire _363;
    wire [131:0] _370;
    wire [63:0] _371;
    wire _299 = 1'b0;
    wire _298 = 1'b0;
    wire _301;
    wire _7;
    reg PHASE_1;
    wire [63:0] _383;
    wire [11:0] address_11;
    wire write_enable_11;
    wire [11:0] address_12;
    wire _570;
    wire read_enable_9;
    wire _568;
    wire write_enable_12;
    wire _572;
    wire [131:0] _577;
    wire [63:0] _578;
    wire [11:0] _563 = 12'b000000000000;
    wire [11:0] address_13;
    wire _561;
    wire write_enable_13;
    wire [63:0] _486;
    wire [63:0] _485;
    wire [63:0] _487;
    wire [63:0] _483;
    wire [63:0] _482;
    wire [63:0] q1_0;
    wire [63:0] _488;
    wire [11:0] address_14;
    wire write_enable_14 = 1'b0;
    wire _473;
    wire read_enable_10;
    wire [11:0] address_15;
    wire _469;
    wire read_enable_11;
    wire _467;
    wire write_enable_15;
    wire _471;
    wire [131:0] _478;
    wire [63:0] _479;
    wire [63:0] data_11 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_12;
    wire [11:0] _461 = 12'b000000000000;
    wire _459;
    wire _458;
    wire _457;
    wire _456;
    wire _455;
    wire _454;
    wire _453;
    wire _452;
    wire _451;
    wire _450;
    wire _449;
    wire _448;
    wire [11:0] _460;
    wire [11:0] address_16;
    wire write_enable_16 = 1'b0;
    wire _445;
    wire read_enable_12;
    wire [63:0] data_13;
    wire [63:0] data_14;
    wire _442;
    wire _441;
    wire _440;
    wire _439;
    wire _438;
    wire _437;
    wire _436;
    wire _435;
    wire _434;
    wire _433;
    wire _432;
    wire _431;
    wire [11:0] _443;
    wire [11:0] address_17;
    wire _428;
    wire read_enable_13;
    wire _426;
    wire write_enable_17;
    wire _430;
    wire [131:0] _465;
    wire [63:0] _466;
    wire _385 = 1'b0;
    wire _384 = 1'b0;
    wire _387;
    wire _11;
    reg PHASE_2;
    wire [63:0] _480;
    wire [11:0] address_18;
    wire _418;
    wire read_enable_14;
    wire write_enable_18;
    wire _420;
    wire [11:0] address_19;
    wire _413;
    wire read_enable_15;
    wire _411;
    wire write_enable_19;
    wire _415;
    wire [131:0] _423;
    wire [63:0] _424;
    wire [63:0] _491;
    wire [63:0] data_15;
    wire [63:0] data_16;
    wire [63:0] data_17;
    wire [63:0] data_18;
    wire [11:0] address_20;
    wire _404;
    wire read_enable_16;
    wire _401;
    wire _402;
    wire write_enable_20;
    wire _406;
    wire [11:0] address_21;
    wire _397;
    wire read_enable_17;
    wire _394;
    wire _395;
    wire write_enable_21;
    wire _399;
    wire [131:0] _409;
    wire [63:0] _410;
    wire _392 = 1'b0;
    wire _391 = 1'b0;
    wire _492;
    wire _13;
    reg PHASE_3;
    wire [63:0] q0_0;
    wire _389 = 1'b0;
    wire _388 = 1'b0;
    reg _390;
    wire [63:0] _481;
    wire [191:0] _490;
    wire [63:0] _493;
    wire [63:0] data_19;
    wire [63:0] data_20;
    wire [63:0] data_21;
    wire [63:0] data_22;
    wire [11:0] address_22;
    wire _557;
    wire _556;
    wire read_enable_18;
    wire _550 = 1'b0;
    wire _549 = 1'b0;
    wire _547 = 1'b0;
    wire _546 = 1'b0;
    wire _544 = 1'b0;
    wire _543 = 1'b0;
    wire _541 = 1'b0;
    wire _540 = 1'b0;
    wire _538 = 1'b0;
    wire _537 = 1'b0;
    wire _535 = 1'b0;
    wire _534 = 1'b0;
    wire _532 = 1'b0;
    wire _531 = 1'b0;
    wire _529 = 1'b0;
    wire _528 = 1'b0;
    wire _526 = 1'b0;
    wire _525 = 1'b0;
    reg _527;
    reg _530;
    reg _533;
    reg _536;
    reg _539;
    reg _542;
    reg _545;
    reg _548;
    reg _551;
    wire _552;
    wire _523 = 1'b0;
    wire _522 = 1'b0;
    wire _520 = 1'b0;
    wire _519 = 1'b0;
    wire _517 = 1'b0;
    wire _516 = 1'b0;
    wire _514 = 1'b0;
    wire _513 = 1'b0;
    wire _511 = 1'b0;
    wire _510 = 1'b0;
    wire _508 = 1'b0;
    wire _507 = 1'b0;
    wire _505 = 1'b0;
    wire _504 = 1'b0;
    wire _502 = 1'b0;
    wire _501 = 1'b0;
    wire _499 = 1'b0;
    wire _498 = 1'b0;
    reg _500;
    reg _503;
    reg _506;
    reg _509;
    reg _512;
    reg _515;
    reg _518;
    reg _521;
    reg _524;
    wire _553;
    wire _554;
    wire write_enable_22;
    wire _559;
    wire [131:0] _566;
    wire [63:0] _567;
    wire _495 = 1'b0;
    wire _494 = 1'b0;
    wire _497;
    wire _15;
    reg PHASE_4;
    wire [63:0] _579;
    wire [11:0] address_23;
    wire write_enable_23;
    wire [11:0] address_24;
    wire _766;
    wire read_enable_19;
    wire _764;
    wire write_enable_24;
    wire _768;
    wire [131:0] _773;
    wire [63:0] _774;
    wire [11:0] _759 = 12'b000000000000;
    wire [11:0] address_25;
    wire _757;
    wire write_enable_25;
    wire [63:0] _682;
    wire [63:0] _681;
    wire [63:0] _683;
    wire [63:0] _679;
    wire [63:0] _678;
    wire [63:0] q1_1;
    wire [63:0] _684;
    wire [11:0] address_26;
    wire write_enable_26 = 1'b0;
    wire _669;
    wire read_enable_20;
    wire [11:0] address_27;
    wire _665;
    wire read_enable_21;
    wire _663;
    wire write_enable_27;
    wire _667;
    wire [131:0] _674;
    wire [63:0] _675;
    wire [63:0] data_23 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_24;
    wire [11:0] _657 = 12'b000000000000;
    wire _655;
    wire _654;
    wire _653;
    wire _652;
    wire _651;
    wire _650;
    wire _649;
    wire _648;
    wire _647;
    wire _646;
    wire _645;
    wire _644;
    wire [11:0] _656;
    wire [11:0] address_28;
    wire write_enable_28 = 1'b0;
    wire _641;
    wire read_enable_22;
    wire [63:0] data_25;
    wire [63:0] data_26;
    wire _638;
    wire _637;
    wire _636;
    wire _635;
    wire _634;
    wire _633;
    wire _632;
    wire _631;
    wire _630;
    wire _629;
    wire _628;
    wire _627;
    wire [11:0] _639;
    wire [11:0] address_29;
    wire _624;
    wire read_enable_23;
    wire _622;
    wire write_enable_29;
    wire _626;
    wire [131:0] _661;
    wire [63:0] _662;
    wire _581 = 1'b0;
    wire _580 = 1'b0;
    wire _583;
    wire _19;
    reg PHASE_5;
    wire [63:0] _676;
    wire [11:0] address_30;
    wire _614;
    wire read_enable_24;
    wire write_enable_30;
    wire _616;
    wire [11:0] address_31;
    wire _609;
    wire read_enable_25;
    wire _607;
    wire write_enable_31;
    wire _611;
    wire [131:0] _619;
    wire [63:0] _620;
    wire [63:0] _687;
    wire [63:0] data_27;
    wire [63:0] data_28;
    wire [63:0] data_29;
    wire [63:0] data_30;
    wire [11:0] address_32;
    wire _600;
    wire read_enable_26;
    wire _597;
    wire _598;
    wire write_enable_32;
    wire _602;
    wire [11:0] address_33;
    wire _593;
    wire read_enable_27;
    wire _590;
    wire _591;
    wire write_enable_33;
    wire _595;
    wire [131:0] _605;
    wire [63:0] _606;
    wire _588 = 1'b0;
    wire _587 = 1'b0;
    wire _688;
    wire _21;
    reg PHASE_6;
    wire [63:0] q0_1;
    wire _585 = 1'b0;
    wire _584 = 1'b0;
    reg _586;
    wire [63:0] _677;
    wire [191:0] _686;
    wire [63:0] _689;
    wire [63:0] data_31;
    wire [63:0] data_32;
    wire [63:0] data_33;
    wire [63:0] data_34;
    wire [11:0] address_34;
    wire _753;
    wire _752;
    wire read_enable_28;
    wire _746 = 1'b0;
    wire _745 = 1'b0;
    wire _743 = 1'b0;
    wire _742 = 1'b0;
    wire _740 = 1'b0;
    wire _739 = 1'b0;
    wire _737 = 1'b0;
    wire _736 = 1'b0;
    wire _734 = 1'b0;
    wire _733 = 1'b0;
    wire _731 = 1'b0;
    wire _730 = 1'b0;
    wire _728 = 1'b0;
    wire _727 = 1'b0;
    wire _725 = 1'b0;
    wire _724 = 1'b0;
    wire _722 = 1'b0;
    wire _721 = 1'b0;
    reg _723;
    reg _726;
    reg _729;
    reg _732;
    reg _735;
    reg _738;
    reg _741;
    reg _744;
    reg _747;
    wire _748;
    wire _719 = 1'b0;
    wire _718 = 1'b0;
    wire _716 = 1'b0;
    wire _715 = 1'b0;
    wire _713 = 1'b0;
    wire _712 = 1'b0;
    wire _710 = 1'b0;
    wire _709 = 1'b0;
    wire _707 = 1'b0;
    wire _706 = 1'b0;
    wire _704 = 1'b0;
    wire _703 = 1'b0;
    wire _701 = 1'b0;
    wire _700 = 1'b0;
    wire _698 = 1'b0;
    wire _697 = 1'b0;
    wire _695 = 1'b0;
    wire _694 = 1'b0;
    reg _696;
    reg _699;
    reg _702;
    reg _705;
    reg _708;
    reg _711;
    reg _714;
    reg _717;
    reg _720;
    wire _749;
    wire _750;
    wire write_enable_34;
    wire _755;
    wire [131:0] _762;
    wire [63:0] _763;
    wire _691 = 1'b0;
    wire _690 = 1'b0;
    wire _693;
    wire _23;
    reg PHASE_7;
    wire [63:0] _775;
    wire [11:0] address_35;
    wire write_enable_35;
    wire [11:0] address_36;
    wire _962;
    wire read_enable_29;
    wire _960;
    wire write_enable_36;
    wire _964;
    wire [131:0] _969;
    wire [63:0] _970;
    wire [11:0] _955 = 12'b000000000000;
    wire [11:0] address_37;
    wire _953;
    wire write_enable_37;
    wire [63:0] _878;
    wire [63:0] _877;
    wire [63:0] _879;
    wire [63:0] _875;
    wire [63:0] _874;
    wire [63:0] q1_2;
    wire [63:0] _880;
    wire [11:0] address_38;
    wire write_enable_38 = 1'b0;
    wire _865;
    wire read_enable_30;
    wire [11:0] address_39;
    wire _861;
    wire read_enable_31;
    wire _859;
    wire write_enable_39;
    wire _863;
    wire [131:0] _870;
    wire [63:0] _871;
    wire [63:0] data_35 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_36;
    wire [11:0] _853 = 12'b000000000000;
    wire _851;
    wire _850;
    wire _849;
    wire _848;
    wire _847;
    wire _846;
    wire _845;
    wire _844;
    wire _843;
    wire _842;
    wire _841;
    wire _840;
    wire [11:0] _852;
    wire [11:0] address_40;
    wire write_enable_40 = 1'b0;
    wire _837;
    wire read_enable_32;
    wire [63:0] data_37;
    wire [63:0] data_38;
    wire _834;
    wire _833;
    wire _832;
    wire _831;
    wire _830;
    wire _829;
    wire _828;
    wire _827;
    wire _826;
    wire _825;
    wire _824;
    wire _823;
    wire [11:0] _835;
    wire [11:0] address_41;
    wire _820;
    wire read_enable_33;
    wire _818;
    wire write_enable_41;
    wire _822;
    wire [131:0] _857;
    wire [63:0] _858;
    wire _777 = 1'b0;
    wire _776 = 1'b0;
    wire _779;
    wire _27;
    reg PHASE_8;
    wire [63:0] _872;
    wire [11:0] address_42;
    wire _810;
    wire read_enable_34;
    wire write_enable_42;
    wire _812;
    wire [11:0] address_43;
    wire _805;
    wire read_enable_35;
    wire _803;
    wire write_enable_43;
    wire _807;
    wire [131:0] _815;
    wire [63:0] _816;
    wire [63:0] _883;
    wire [63:0] data_39;
    wire [63:0] data_40;
    wire [63:0] data_41;
    wire [63:0] data_42;
    wire [11:0] address_44;
    wire _796;
    wire read_enable_36;
    wire _793;
    wire _794;
    wire write_enable_44;
    wire _798;
    wire [11:0] address_45;
    wire _789;
    wire read_enable_37;
    wire _786;
    wire _787;
    wire write_enable_45;
    wire _791;
    wire [131:0] _801;
    wire [63:0] _802;
    wire _784 = 1'b0;
    wire _783 = 1'b0;
    wire _884;
    wire _29;
    reg PHASE_9;
    wire [63:0] q0_2;
    wire _781 = 1'b0;
    wire _780 = 1'b0;
    reg _782;
    wire [63:0] _873;
    wire [191:0] _882;
    wire [63:0] _885;
    wire [63:0] data_43;
    wire [63:0] data_44;
    wire [63:0] data_45;
    wire [63:0] data_46;
    wire [11:0] address_46;
    wire _949;
    wire _948;
    wire read_enable_38;
    wire _942 = 1'b0;
    wire _941 = 1'b0;
    wire _939 = 1'b0;
    wire _938 = 1'b0;
    wire _936 = 1'b0;
    wire _935 = 1'b0;
    wire _933 = 1'b0;
    wire _932 = 1'b0;
    wire _930 = 1'b0;
    wire _929 = 1'b0;
    wire _927 = 1'b0;
    wire _926 = 1'b0;
    wire _924 = 1'b0;
    wire _923 = 1'b0;
    wire _921 = 1'b0;
    wire _920 = 1'b0;
    wire _918 = 1'b0;
    wire _917 = 1'b0;
    reg _919;
    reg _922;
    reg _925;
    reg _928;
    reg _931;
    reg _934;
    reg _937;
    reg _940;
    reg _943;
    wire _944;
    wire _915 = 1'b0;
    wire _914 = 1'b0;
    wire _912 = 1'b0;
    wire _911 = 1'b0;
    wire _909 = 1'b0;
    wire _908 = 1'b0;
    wire _906 = 1'b0;
    wire _905 = 1'b0;
    wire _903 = 1'b0;
    wire _902 = 1'b0;
    wire _900 = 1'b0;
    wire _899 = 1'b0;
    wire _897 = 1'b0;
    wire _896 = 1'b0;
    wire _894 = 1'b0;
    wire _893 = 1'b0;
    wire _891 = 1'b0;
    wire _890 = 1'b0;
    reg _892;
    reg _895;
    reg _898;
    reg _901;
    reg _904;
    reg _907;
    reg _910;
    reg _913;
    reg _916;
    wire _945;
    wire _946;
    wire write_enable_46;
    wire _951;
    wire [131:0] _958;
    wire [63:0] _959;
    wire _887 = 1'b0;
    wire _886 = 1'b0;
    wire _889;
    wire _31;
    reg PHASE_10;
    wire [63:0] _971;
    wire [11:0] address_47;
    wire write_enable_47;
    wire [11:0] address_48;
    wire _1158;
    wire read_enable_39;
    wire _1156;
    wire write_enable_48;
    wire _1160;
    wire [131:0] _1165;
    wire [63:0] _1166;
    wire [11:0] _1151 = 12'b000000000000;
    wire [11:0] address_49;
    wire _1149;
    wire write_enable_49;
    wire [63:0] _1074;
    wire [63:0] _1073;
    wire [63:0] _1075;
    wire [63:0] _1071;
    wire [63:0] _1070;
    wire [63:0] q1_3;
    wire [63:0] _1076;
    wire [11:0] address_50;
    wire write_enable_50 = 1'b0;
    wire _1061;
    wire read_enable_40;
    wire [11:0] address_51;
    wire _1057;
    wire read_enable_41;
    wire _1055;
    wire write_enable_51;
    wire _1059;
    wire [131:0] _1066;
    wire [63:0] _1067;
    wire [63:0] data_47 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_48;
    wire [11:0] _1049 = 12'b000000000000;
    wire _1047;
    wire _1046;
    wire _1045;
    wire _1044;
    wire _1043;
    wire _1042;
    wire _1041;
    wire _1040;
    wire _1039;
    wire _1038;
    wire _1037;
    wire _1036;
    wire [11:0] _1048;
    wire [11:0] address_52;
    wire write_enable_52 = 1'b0;
    wire _1033;
    wire read_enable_42;
    wire [63:0] data_49;
    wire [63:0] data_50;
    wire _1030;
    wire _1029;
    wire _1028;
    wire _1027;
    wire _1026;
    wire _1025;
    wire _1024;
    wire _1023;
    wire _1022;
    wire _1021;
    wire _1020;
    wire _1019;
    wire [11:0] _1031;
    wire [11:0] address_53;
    wire _1016;
    wire read_enable_43;
    wire _1014;
    wire write_enable_53;
    wire _1018;
    wire [131:0] _1053;
    wire [63:0] _1054;
    wire _973 = 1'b0;
    wire _972 = 1'b0;
    wire _975;
    wire _35;
    reg PHASE_11;
    wire [63:0] _1068;
    wire [11:0] address_54;
    wire _1006;
    wire read_enable_44;
    wire write_enable_54;
    wire _1008;
    wire [11:0] address_55;
    wire _1001;
    wire read_enable_45;
    wire _999;
    wire write_enable_55;
    wire _1003;
    wire [131:0] _1011;
    wire [63:0] _1012;
    wire [63:0] _1079;
    wire [63:0] data_51;
    wire [63:0] data_52;
    wire [63:0] data_53;
    wire [63:0] data_54;
    wire [11:0] address_56;
    wire _992;
    wire read_enable_46;
    wire _989;
    wire _990;
    wire write_enable_56;
    wire _994;
    wire [11:0] address_57;
    wire _985;
    wire read_enable_47;
    wire _982;
    wire _983;
    wire write_enable_57;
    wire _987;
    wire [131:0] _997;
    wire [63:0] _998;
    wire _980 = 1'b0;
    wire _979 = 1'b0;
    wire _1080;
    wire _37;
    reg PHASE_12;
    wire [63:0] q0_3;
    wire _977 = 1'b0;
    wire _976 = 1'b0;
    reg _978;
    wire [63:0] _1069;
    wire [191:0] _1078;
    wire [63:0] _1081;
    wire [63:0] data_55;
    wire [63:0] data_56;
    wire [63:0] data_57;
    wire [63:0] data_58;
    wire [11:0] address_58;
    wire _1145;
    wire _1144;
    wire read_enable_48;
    wire _1138 = 1'b0;
    wire _1137 = 1'b0;
    wire _1135 = 1'b0;
    wire _1134 = 1'b0;
    wire _1132 = 1'b0;
    wire _1131 = 1'b0;
    wire _1129 = 1'b0;
    wire _1128 = 1'b0;
    wire _1126 = 1'b0;
    wire _1125 = 1'b0;
    wire _1123 = 1'b0;
    wire _1122 = 1'b0;
    wire _1120 = 1'b0;
    wire _1119 = 1'b0;
    wire _1117 = 1'b0;
    wire _1116 = 1'b0;
    wire _1114 = 1'b0;
    wire _1113 = 1'b0;
    reg _1115;
    reg _1118;
    reg _1121;
    reg _1124;
    reg _1127;
    reg _1130;
    reg _1133;
    reg _1136;
    reg _1139;
    wire _1140;
    wire _1111 = 1'b0;
    wire _1110 = 1'b0;
    wire _1108 = 1'b0;
    wire _1107 = 1'b0;
    wire _1105 = 1'b0;
    wire _1104 = 1'b0;
    wire _1102 = 1'b0;
    wire _1101 = 1'b0;
    wire _1099 = 1'b0;
    wire _1098 = 1'b0;
    wire _1096 = 1'b0;
    wire _1095 = 1'b0;
    wire _1093 = 1'b0;
    wire _1092 = 1'b0;
    wire _1090 = 1'b0;
    wire _1089 = 1'b0;
    wire _1087 = 1'b0;
    wire _1086 = 1'b0;
    reg _1088;
    reg _1091;
    reg _1094;
    reg _1097;
    reg _1100;
    reg _1103;
    reg _1106;
    reg _1109;
    reg _1112;
    wire _1141;
    wire _1142;
    wire write_enable_58;
    wire _1147;
    wire [131:0] _1154;
    wire [63:0] _1155;
    wire _1083 = 1'b0;
    wire _1082 = 1'b0;
    wire _1085;
    wire _39;
    reg PHASE_13;
    wire [63:0] _1167;
    wire [11:0] address_59;
    wire write_enable_59;
    wire [11:0] address_60;
    wire _1354;
    wire read_enable_49;
    wire _1352;
    wire write_enable_60;
    wire _1356;
    wire [131:0] _1361;
    wire [63:0] _1362;
    wire [11:0] _1347 = 12'b000000000000;
    wire [11:0] address_61;
    wire _1345;
    wire write_enable_61;
    wire [63:0] _1270;
    wire [63:0] _1269;
    wire [63:0] _1271;
    wire [63:0] _1267;
    wire [63:0] _1266;
    wire [63:0] q1_4;
    wire [63:0] _1272;
    wire [11:0] address_62;
    wire write_enable_62 = 1'b0;
    wire _1257;
    wire read_enable_50;
    wire [11:0] address_63;
    wire _1253;
    wire read_enable_51;
    wire _1251;
    wire write_enable_63;
    wire _1255;
    wire [131:0] _1262;
    wire [63:0] _1263;
    wire [63:0] data_59 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_60;
    wire [11:0] _1245 = 12'b000000000000;
    wire _1243;
    wire _1242;
    wire _1241;
    wire _1240;
    wire _1239;
    wire _1238;
    wire _1237;
    wire _1236;
    wire _1235;
    wire _1234;
    wire _1233;
    wire _1232;
    wire [11:0] _1244;
    wire [11:0] address_64;
    wire write_enable_64 = 1'b0;
    wire _1229;
    wire read_enable_52;
    wire [63:0] data_61;
    wire [63:0] data_62;
    wire _1226;
    wire _1225;
    wire _1224;
    wire _1223;
    wire _1222;
    wire _1221;
    wire _1220;
    wire _1219;
    wire _1218;
    wire _1217;
    wire _1216;
    wire _1215;
    wire [11:0] _1227;
    wire [11:0] address_65;
    wire _1212;
    wire read_enable_53;
    wire _1210;
    wire write_enable_65;
    wire _1214;
    wire [131:0] _1249;
    wire [63:0] _1250;
    wire _1169 = 1'b0;
    wire _1168 = 1'b0;
    wire _1171;
    wire _43;
    reg PHASE_14;
    wire [63:0] _1264;
    wire [11:0] address_66;
    wire _1202;
    wire read_enable_54;
    wire write_enable_66;
    wire _1204;
    wire [11:0] address_67;
    wire _1197;
    wire read_enable_55;
    wire _1195;
    wire write_enable_67;
    wire _1199;
    wire [131:0] _1207;
    wire [63:0] _1208;
    wire [63:0] _1275;
    wire [63:0] data_63;
    wire [63:0] data_64;
    wire [63:0] data_65;
    wire [63:0] data_66;
    wire [11:0] address_68;
    wire _1188;
    wire read_enable_56;
    wire _1185;
    wire _1186;
    wire write_enable_68;
    wire _1190;
    wire [11:0] address_69;
    wire _1181;
    wire read_enable_57;
    wire _1178;
    wire _1179;
    wire write_enable_69;
    wire _1183;
    wire [131:0] _1193;
    wire [63:0] _1194;
    wire _1176 = 1'b0;
    wire _1175 = 1'b0;
    wire _1276;
    wire _45;
    reg PHASE_15;
    wire [63:0] q0_4;
    wire _1173 = 1'b0;
    wire _1172 = 1'b0;
    reg _1174;
    wire [63:0] _1265;
    wire [191:0] _1274;
    wire [63:0] _1277;
    wire [63:0] data_67;
    wire [63:0] data_68;
    wire [63:0] data_69;
    wire [63:0] data_70;
    wire [11:0] address_70;
    wire _1341;
    wire _1340;
    wire read_enable_58;
    wire _1334 = 1'b0;
    wire _1333 = 1'b0;
    wire _1331 = 1'b0;
    wire _1330 = 1'b0;
    wire _1328 = 1'b0;
    wire _1327 = 1'b0;
    wire _1325 = 1'b0;
    wire _1324 = 1'b0;
    wire _1322 = 1'b0;
    wire _1321 = 1'b0;
    wire _1319 = 1'b0;
    wire _1318 = 1'b0;
    wire _1316 = 1'b0;
    wire _1315 = 1'b0;
    wire _1313 = 1'b0;
    wire _1312 = 1'b0;
    wire _1310 = 1'b0;
    wire _1309 = 1'b0;
    reg _1311;
    reg _1314;
    reg _1317;
    reg _1320;
    reg _1323;
    reg _1326;
    reg _1329;
    reg _1332;
    reg _1335;
    wire _1336;
    wire _1307 = 1'b0;
    wire _1306 = 1'b0;
    wire _1304 = 1'b0;
    wire _1303 = 1'b0;
    wire _1301 = 1'b0;
    wire _1300 = 1'b0;
    wire _1298 = 1'b0;
    wire _1297 = 1'b0;
    wire _1295 = 1'b0;
    wire _1294 = 1'b0;
    wire _1292 = 1'b0;
    wire _1291 = 1'b0;
    wire _1289 = 1'b0;
    wire _1288 = 1'b0;
    wire _1286 = 1'b0;
    wire _1285 = 1'b0;
    wire _1283 = 1'b0;
    wire _1282 = 1'b0;
    reg _1284;
    reg _1287;
    reg _1290;
    reg _1293;
    reg _1296;
    reg _1299;
    reg _1302;
    reg _1305;
    reg _1308;
    wire _1337;
    wire _1338;
    wire write_enable_70;
    wire _1343;
    wire [131:0] _1350;
    wire [63:0] _1351;
    wire _1279 = 1'b0;
    wire _1278 = 1'b0;
    wire _1281;
    wire _47;
    reg PHASE_16;
    wire [63:0] _1363;
    wire [11:0] address_71;
    wire write_enable_71;
    wire [11:0] address_72;
    wire _1550;
    wire read_enable_59;
    wire _1548;
    wire write_enable_72;
    wire _1552;
    wire [131:0] _1557;
    wire [63:0] _1558;
    wire [11:0] _1543 = 12'b000000000000;
    wire [11:0] address_73;
    wire _1541;
    wire write_enable_73;
    wire [63:0] _1466;
    wire [63:0] _1465;
    wire [63:0] _1467;
    wire [63:0] _1463;
    wire [63:0] _1462;
    wire [63:0] q1_5;
    wire [63:0] _1468;
    wire [11:0] address_74;
    wire write_enable_74 = 1'b0;
    wire _1453;
    wire read_enable_60;
    wire [11:0] address_75;
    wire _1449;
    wire read_enable_61;
    wire _1447;
    wire write_enable_75;
    wire _1451;
    wire [131:0] _1458;
    wire [63:0] _1459;
    wire [63:0] data_71 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_72;
    wire [11:0] _1441 = 12'b000000000000;
    wire _1439;
    wire _1438;
    wire _1437;
    wire _1436;
    wire _1435;
    wire _1434;
    wire _1433;
    wire _1432;
    wire _1431;
    wire _1430;
    wire _1429;
    wire _1428;
    wire [11:0] _1440;
    wire [11:0] address_76;
    wire write_enable_76 = 1'b0;
    wire _1425;
    wire read_enable_62;
    wire [63:0] data_73;
    wire [63:0] data_74;
    wire _1422;
    wire _1421;
    wire _1420;
    wire _1419;
    wire _1418;
    wire _1417;
    wire _1416;
    wire _1415;
    wire _1414;
    wire _1413;
    wire _1412;
    wire _1411;
    wire [11:0] _1423;
    wire [11:0] address_77;
    wire _1408;
    wire read_enable_63;
    wire _1406;
    wire write_enable_77;
    wire _1410;
    wire [131:0] _1445;
    wire [63:0] _1446;
    wire _1365 = 1'b0;
    wire _1364 = 1'b0;
    wire _1367;
    wire _51;
    reg PHASE_17;
    wire [63:0] _1460;
    wire [11:0] address_78;
    wire _1398;
    wire read_enable_64;
    wire write_enable_78;
    wire _1400;
    wire [11:0] address_79;
    wire _1393;
    wire read_enable_65;
    wire _1391;
    wire write_enable_79;
    wire _1395;
    wire [131:0] _1403;
    wire [63:0] _1404;
    wire [63:0] _1471;
    wire [63:0] data_75;
    wire [63:0] data_76;
    wire [63:0] data_77;
    wire [63:0] data_78;
    wire [11:0] address_80;
    wire _1384;
    wire read_enable_66;
    wire _1381;
    wire _1382;
    wire write_enable_80;
    wire _1386;
    wire [11:0] address_81;
    wire _1377;
    wire read_enable_67;
    wire _1374;
    wire _1375;
    wire write_enable_81;
    wire _1379;
    wire [131:0] _1389;
    wire [63:0] _1390;
    wire _1372 = 1'b0;
    wire _1371 = 1'b0;
    wire _1472;
    wire _53;
    reg PHASE_18;
    wire [63:0] q0_5;
    wire _1369 = 1'b0;
    wire _1368 = 1'b0;
    reg _1370;
    wire [63:0] _1461;
    wire [191:0] _1470;
    wire [63:0] _1473;
    wire [63:0] data_79;
    wire [63:0] data_80;
    wire [63:0] data_81;
    wire [63:0] data_82;
    wire [11:0] address_82;
    wire _1537;
    wire _1536;
    wire read_enable_68;
    wire _1530 = 1'b0;
    wire _1529 = 1'b0;
    wire _1527 = 1'b0;
    wire _1526 = 1'b0;
    wire _1524 = 1'b0;
    wire _1523 = 1'b0;
    wire _1521 = 1'b0;
    wire _1520 = 1'b0;
    wire _1518 = 1'b0;
    wire _1517 = 1'b0;
    wire _1515 = 1'b0;
    wire _1514 = 1'b0;
    wire _1512 = 1'b0;
    wire _1511 = 1'b0;
    wire _1509 = 1'b0;
    wire _1508 = 1'b0;
    wire _1506 = 1'b0;
    wire _1505 = 1'b0;
    reg _1507;
    reg _1510;
    reg _1513;
    reg _1516;
    reg _1519;
    reg _1522;
    reg _1525;
    reg _1528;
    reg _1531;
    wire _1532;
    wire _1503 = 1'b0;
    wire _1502 = 1'b0;
    wire _1500 = 1'b0;
    wire _1499 = 1'b0;
    wire _1497 = 1'b0;
    wire _1496 = 1'b0;
    wire _1494 = 1'b0;
    wire _1493 = 1'b0;
    wire _1491 = 1'b0;
    wire _1490 = 1'b0;
    wire _1488 = 1'b0;
    wire _1487 = 1'b0;
    wire _1485 = 1'b0;
    wire _1484 = 1'b0;
    wire _1482 = 1'b0;
    wire _1481 = 1'b0;
    wire _1479 = 1'b0;
    wire _1478 = 1'b0;
    reg _1480;
    reg _1483;
    reg _1486;
    reg _1489;
    reg _1492;
    reg _1495;
    reg _1498;
    reg _1501;
    reg _1504;
    wire _1533;
    wire _1534;
    wire write_enable_82;
    wire _1539;
    wire [131:0] _1546;
    wire [63:0] _1547;
    wire _1475 = 1'b0;
    wire _1474 = 1'b0;
    wire _1477;
    wire _55;
    reg PHASE_19;
    wire [63:0] _1559;
    wire [11:0] address_83;
    wire write_enable_83;
    wire [11:0] address_84;
    wire _1746;
    wire read_enable_69;
    wire _1744;
    wire write_enable_84;
    wire _1748;
    wire [131:0] _1753;
    wire [63:0] _1754;
    wire [11:0] _1739 = 12'b000000000000;
    wire [11:0] address_85;
    wire _1737;
    wire write_enable_85;
    wire [3:0] _292;
    wire _291;
    wire _289;
    wire [63:0] _288;
    wire [63:0] _287;
    wire [63:0] _286;
    wire [63:0] _285;
    wire [63:0] _284;
    wire [63:0] _283;
    wire [63:0] _282;
    wire [63:0] _1662;
    wire [63:0] _1661;
    wire [63:0] _1663;
    wire [63:0] _1659;
    wire [63:0] _1658;
    wire [63:0] q1_6;
    wire [63:0] _1664;
    wire [11:0] address_86;
    wire write_enable_86 = 1'b0;
    wire _1649;
    wire read_enable_70;
    wire [11:0] address_87;
    wire _1645;
    wire read_enable_71;
    wire _1643;
    wire write_enable_87;
    wire _1647;
    wire [131:0] _1654;
    wire [63:0] _1655;
    wire [63:0] data_83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_84;
    wire [11:0] _1637 = 12'b000000000000;
    wire _1635;
    wire _1634;
    wire _1633;
    wire _1632;
    wire _1631;
    wire _1630;
    wire _1629;
    wire _1628;
    wire _1627;
    wire _1626;
    wire _1625;
    wire _1624;
    wire [11:0] _1636;
    wire [11:0] address_88;
    wire write_enable_88 = 1'b0;
    wire _1621;
    wire read_enable_72;
    wire [63:0] data_85;
    wire [63:0] data_86;
    wire [11:0] _60;
    wire _1618;
    wire _1617;
    wire _1616;
    wire _1615;
    wire _1614;
    wire _1613;
    wire _1612;
    wire _1611;
    wire _1610;
    wire _1609;
    wire _1608;
    wire _1607;
    wire [11:0] _1619;
    wire [11:0] address_89;
    wire _1604;
    wire read_enable_73;
    wire [7:0] _62;
    wire _1602;
    wire write_enable_89;
    wire _1606;
    wire [131:0] _1641;
    wire [63:0] _1642;
    wire _1561 = 1'b0;
    wire _1560 = 1'b0;
    wire _1563;
    wire _63;
    reg PHASE_20;
    wire [63:0] _1656;
    wire [11:0] address_90;
    wire _1594;
    wire read_enable_74;
    wire write_enable_90;
    wire _1596;
    wire [11:0] address_91;
    wire _1589;
    wire read_enable_75;
    wire _1587;
    wire write_enable_91;
    wire _1591;
    wire [131:0] _1599;
    wire [63:0] _1600;
    wire [63:0] _1667;
    wire [63:0] data_87;
    wire [63:0] data_88;
    wire [63:0] data_89;
    wire [63:0] data_90;
    wire [11:0] _198 = 12'b000000000000;
    wire [11:0] _197 = 12'b000000000000;
    wire [11:0] _195 = 12'b000000000000;
    wire [11:0] _194 = 12'b000000000000;
    wire [11:0] _192 = 12'b000000000000;
    wire [11:0] _191 = 12'b000000000000;
    wire [11:0] _189 = 12'b000000000000;
    wire [11:0] _188 = 12'b000000000000;
    wire [11:0] _186 = 12'b000000000000;
    wire [11:0] _185 = 12'b000000000000;
    wire [11:0] _183 = 12'b000000000000;
    wire [11:0] _182 = 12'b000000000000;
    wire [11:0] _180 = 12'b000000000000;
    wire [11:0] _179 = 12'b000000000000;
    wire [11:0] _177 = 12'b000000000000;
    wire [11:0] _176 = 12'b000000000000;
    wire [11:0] _174 = 12'b000000000000;
    wire [11:0] _173 = 12'b000000000000;
    reg [11:0] _175;
    reg [11:0] _178;
    reg [11:0] _181;
    reg [11:0] _184;
    reg [11:0] _187;
    reg [11:0] _190;
    reg [11:0] _193;
    reg [11:0] _196;
    reg [11:0] _199;
    wire [11:0] _172;
    wire [11:0] address_92;
    wire _1580;
    wire read_enable_76;
    wire _1577;
    wire _1578;
    wire write_enable_92;
    wire _1582;
    wire [11:0] address_93;
    wire _1573;
    wire read_enable_77;
    wire _1570;
    wire _1571;
    wire write_enable_93;
    wire _1575;
    wire [131:0] _1585;
    wire [63:0] _1586;
    wire _99;
    wire _1568 = 1'b0;
    wire _1567 = 1'b0;
    wire _1668;
    wire _65;
    reg PHASE_21;
    wire [63:0] q0_6;
    wire _1565 = 1'b0;
    wire _1564 = 1'b0;
    wire _92;
    reg _1566;
    wire [63:0] _1657;
    wire [191:0] _1666;
    wire [63:0] _1669;
    wire [63:0] data_91;
    wire [63:0] data_92;
    wire [63:0] data_93;
    wire [63:0] data_94;
    wire [11:0] _163 = 12'b000000000000;
    wire [11:0] _162 = 12'b000000000000;
    wire [11:0] _160 = 12'b000000000000;
    wire [11:0] _159 = 12'b000000000000;
    wire [11:0] _157 = 12'b000000000000;
    wire [11:0] _156 = 12'b000000000000;
    wire [11:0] _154 = 12'b000000000000;
    wire [11:0] _153 = 12'b000000000000;
    wire [11:0] _151 = 12'b000000000000;
    wire [11:0] _150 = 12'b000000000000;
    wire [11:0] _148 = 12'b000000000000;
    wire [11:0] _147 = 12'b000000000000;
    wire [11:0] _145 = 12'b000000000000;
    wire [11:0] _144 = 12'b000000000000;
    wire [11:0] _142 = 12'b000000000000;
    wire [11:0] _141 = 12'b000000000000;
    wire [11:0] _139 = 12'b000000000000;
    wire [11:0] _138 = 12'b000000000000;
    wire [11:0] _137;
    reg [11:0] _140;
    reg [11:0] _143;
    reg [11:0] _146;
    reg [11:0] _149;
    reg [11:0] _152;
    reg [11:0] _155;
    reg [11:0] _158;
    reg [11:0] _161;
    reg [11:0] _164;
    wire [11:0] _68;
    wire [11:0] address_94;
    wire _1733;
    wire [7:0] _70;
    wire _1732;
    wire read_enable_78;
    wire _1726 = 1'b0;
    wire _1725 = 1'b0;
    wire _1723 = 1'b0;
    wire _1722 = 1'b0;
    wire _1720 = 1'b0;
    wire _1719 = 1'b0;
    wire _1717 = 1'b0;
    wire _1716 = 1'b0;
    wire _1714 = 1'b0;
    wire _1713 = 1'b0;
    wire _1711 = 1'b0;
    wire _1710 = 1'b0;
    wire _1708 = 1'b0;
    wire _1707 = 1'b0;
    wire _1705 = 1'b0;
    wire _1704 = 1'b0;
    wire _1702 = 1'b0;
    wire _1701 = 1'b0;
    wire _290;
    reg _1703;
    reg _1706;
    reg _1709;
    reg _1712;
    reg _1715;
    reg _1718;
    reg _1721;
    reg _1724;
    reg _1727;
    wire _1728;
    wire _1699 = 1'b0;
    wire _1698 = 1'b0;
    wire _1696 = 1'b0;
    wire _1695 = 1'b0;
    wire _1693 = 1'b0;
    wire _1692 = 1'b0;
    wire _1690 = 1'b0;
    wire _1689 = 1'b0;
    wire _1687 = 1'b0;
    wire _1686 = 1'b0;
    wire _1684 = 1'b0;
    wire _1683 = 1'b0;
    wire _1681 = 1'b0;
    wire _1680 = 1'b0;
    wire _1678 = 1'b0;
    wire _1677 = 1'b0;
    wire _1675 = 1'b0;
    wire _1674 = 1'b0;
    wire _130;
    reg _1676;
    reg _1679;
    reg _1682;
    reg _1685;
    reg _1688;
    reg _1691;
    reg _1694;
    reg _1697;
    reg _1700;
    wire _1729;
    wire _128 = 1'b0;
    wire _127 = 1'b0;
    wire _125 = 1'b0;
    wire _124 = 1'b0;
    wire _122 = 1'b0;
    wire _121 = 1'b0;
    wire _119 = 1'b0;
    wire _118 = 1'b0;
    wire _116 = 1'b0;
    wire _115 = 1'b0;
    wire _113 = 1'b0;
    wire _112 = 1'b0;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire vdd = 1'b1;
    wire _104 = 1'b0;
    wire _103 = 1'b0;
    wire _102;
    reg _105;
    reg _108;
    reg _111;
    reg _114;
    reg _117;
    reg _120;
    reg _123;
    reg _126;
    reg _129;
    wire _1730;
    wire write_enable_94;
    wire _1735;
    wire gnd = 1'b0;
    wire [131:0] _1742;
    wire [63:0] _1743;
    wire _72;
    wire _1671 = 1'b0;
    wire _1670 = 1'b0;
    wire _1673;
    wire _73;
    reg PHASE_22;
    wire [63:0] _1755;
    wire _76;
    wire _78;
    wire _80;
    wire _82;
    wire _84;
    wire [523:0] _91;
    wire _1756;

    /* logic */
    assign address = _372 ? _199 : _367;
    assign write_enable = _365 & _372;
    assign address_0 = _372 ? _164 : _68;
    assign _374 = ~ _372;
    assign read_enable = _360 & _374;
    assign _372 = ~ PHASE_1;
    assign write_enable_0 = _358 & _372;
    assign _376 = write_enable_0 | read_enable;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_376), .regcea(vdd), .wea(write_enable_0), .addra(address_0), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable), .regceb(vdd), .web(write_enable), .addrb(address), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_381[131:131]), .sbiterrb(_381[130:130]), .doutb(_381[129:66]), .dbiterra(_381[65:65]), .sbiterra(_381[64:64]), .douta(_381[63:0]) );
    assign _382 = _381[63:0];
    assign address_1 = PHASE_1 ? _199 : _367;
    assign _365 = _129 & _328;
    assign write_enable_1 = _365 & PHASE_1;
    assign _279 = _271[129:66];
    assign _278 = _258[129:66];
    assign _280 = PHASE ? _279 : _278;
    assign _276 = _216[129:66];
    assign _275 = _202[129:66];
    assign q1 = PHASE_0 ? _276 : _275;
    assign _281 = _96 ? _280 : q1;
    assign address_2 = _260 ? _254 : _253;
    assign _266 = ~ _260;
    assign read_enable_0 = _102 & _266;
    assign address_3 = _260 ? _60 : _236;
    assign _262 = ~ _260;
    assign read_enable_1 = _102 & _262;
    assign _260 = ~ PHASE;
    assign write_enable_3 = _219 & _260;
    assign _264 = write_enable_3 | read_enable_1;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_0
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_264), .regcea(vdd), .wea(write_enable_3), .addra(address_3), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_0), .regceb(vdd), .web(write_enable_2), .addrb(address_2), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_271[131:131]), .sbiterrb(_271[130:130]), .doutb(_271[129:66]), .dbiterra(_271[65:65]), .sbiterra(_271[64:64]), .douta(_271[63:0]) );
    assign _272 = _271[63:0];
    assign _252 = _172[11:11];
    assign _251 = _172[10:10];
    assign _250 = _172[9:9];
    assign _249 = _172[8:8];
    assign _248 = _172[7:7];
    assign _247 = _172[6:6];
    assign _246 = _172[5:5];
    assign _245 = _172[4:4];
    assign _244 = _172[3:3];
    assign _243 = _172[2:2];
    assign _242 = _172[1:1];
    assign _241 = _172[0:0];
    assign _253 = { _241, _242, _243, _244, _245, _246, _247, _248, _249, _250, _251, _252 };
    assign address_4 = PHASE ? _254 : _253;
    assign _238 = ~ PHASE;
    assign read_enable_2 = _102 & _238;
    assign data_1 = wr_d7;
    assign _235 = _137[11:11];
    assign _234 = _137[10:10];
    assign _233 = _137[9:9];
    assign _232 = _137[8:8];
    assign _231 = _137[7:7];
    assign _230 = _137[6:6];
    assign _229 = _137[5:5];
    assign _228 = _137[4:4];
    assign _227 = _137[3:3];
    assign _226 = _137[2:2];
    assign _225 = _137[1:1];
    assign _224 = _137[0:0];
    assign _236 = { _224, _225, _226, _227, _228, _229, _230, _231, _232, _233, _234, _235 };
    assign address_5 = PHASE ? _60 : _236;
    assign _221 = ~ PHASE;
    assign read_enable_3 = _102 & _221;
    assign _219 = _62[7:7];
    assign write_enable_5 = _219 & PHASE;
    assign _223 = write_enable_5 | read_enable_3;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_1
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_223), .regcea(vdd), .wea(write_enable_5), .addra(address_5), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_2), .regceb(vdd), .web(write_enable_4), .addrb(address_4), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_258[131:131]), .sbiterrb(_258[130:130]), .doutb(_258[129:66]), .dbiterra(_258[65:65]), .sbiterra(_258[64:64]), .douta(_258[63:0]) );
    assign _259 = _258[63:0];
    assign _89 = ~ PHASE;
    assign _3 = _89;
    always @(posedge _84) begin
        if (_82)
            PHASE <= _87;
        else
            if (_72)
                PHASE <= _3;
    end
    assign _273 = PHASE ? _272 : _259;
    assign address_6 = _204 ? _199 : _172;
    assign _211 = ~ _204;
    assign read_enable_4 = _102 & _211;
    assign write_enable_6 = _167 & _204;
    assign _213 = write_enable_6 | read_enable_4;
    assign address_7 = _204 ? _164 : _137;
    assign _206 = ~ _204;
    assign read_enable_5 = _102 & _206;
    assign _204 = ~ PHASE_0;
    assign write_enable_7 = _132 & _204;
    assign _208 = write_enable_7 | read_enable_5;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_2
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_208), .regcea(vdd), .wea(write_enable_7), .addra(address_7), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_213), .regceb(vdd), .web(write_enable_6), .addrb(address_6), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_216[131:131]), .sbiterrb(_216[130:130]), .doutb(_216[129:66]), .dbiterra(_216[65:65]), .sbiterra(_216[64:64]), .douta(_216[63:0]) );
    assign _217 = _216[63:0];
    assign _295 = _294[127:64];
    assign data_3 = _295;
    assign address_8 = PHASE_0 ? _199 : _172;
    assign _169 = ~ PHASE_0;
    assign read_enable_6 = _102 & _169;
    assign _166 = ~ _130;
    assign _167 = _129 & _166;
    assign write_enable_8 = _167 & PHASE_0;
    assign _171 = write_enable_8 | read_enable_6;
    assign address_9 = PHASE_0 ? _164 : _137;
    assign _134 = ~ PHASE_0;
    assign read_enable_7 = _102 & _134;
    assign _131 = ~ _130;
    assign _132 = _129 & _131;
    assign write_enable_9 = _132 & PHASE_0;
    assign _136 = write_enable_9 | read_enable_7;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_3
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_136), .regcea(vdd), .wea(write_enable_9), .addra(address_9), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_171), .regceb(vdd), .web(write_enable_8), .addrb(address_8), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_202[131:131]), .sbiterrb(_202[130:130]), .doutb(_202[129:66]), .dbiterra(_202[65:65]), .sbiterra(_202[64:64]), .douta(_202[63:0]) );
    assign _203 = _202[63:0];
    assign _296 = ~ PHASE_0;
    assign _5 = _296;
    always @(posedge _84) begin
        if (_82)
            PHASE_0 <= _98;
        else
            if (_99)
                PHASE_0 <= _5;
    end
    assign q0 = PHASE_0 ? _217 : _203;
    always @(posedge _84) begin
        if (_82)
            _96 <= _94;
        else
            _96 <= _92;
    end
    assign _274 = _96 ? _273 : q0;
    dp_22
        dp_6
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_274), .d2(_281), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_294[191:128]), .q2(_294[127:64]), .q1(_294[63:0]) );
    assign _297 = _294[63:0];
    assign data_7 = _297;
    assign address_10 = PHASE_1 ? _164 : _68;
    assign _361 = ~ PHASE_1;
    assign _360 = _70[7:7];
    assign read_enable_8 = _360 & _361;
    always @(posedge _84) begin
        if (_82)
            _331 <= _330;
        else
            _331 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _334 <= _333;
        else
            _334 <= _331;
    end
    always @(posedge _84) begin
        if (_82)
            _337 <= _336;
        else
            _337 <= _334;
    end
    always @(posedge _84) begin
        if (_82)
            _340 <= _339;
        else
            _340 <= _337;
    end
    always @(posedge _84) begin
        if (_82)
            _343 <= _342;
        else
            _343 <= _340;
    end
    always @(posedge _84) begin
        if (_82)
            _346 <= _345;
        else
            _346 <= _343;
    end
    always @(posedge _84) begin
        if (_82)
            _349 <= _348;
        else
            _349 <= _346;
    end
    always @(posedge _84) begin
        if (_82)
            _352 <= _351;
        else
            _352 <= _349;
    end
    always @(posedge _84) begin
        if (_82)
            _355 <= _354;
        else
            _355 <= _352;
    end
    assign _356 = ~ _355;
    always @(posedge _84) begin
        if (_82)
            _304 <= _303;
        else
            _304 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _307 <= _306;
        else
            _307 <= _304;
    end
    always @(posedge _84) begin
        if (_82)
            _310 <= _309;
        else
            _310 <= _307;
    end
    always @(posedge _84) begin
        if (_82)
            _313 <= _312;
        else
            _313 <= _310;
    end
    always @(posedge _84) begin
        if (_82)
            _316 <= _315;
        else
            _316 <= _313;
    end
    always @(posedge _84) begin
        if (_82)
            _319 <= _318;
        else
            _319 <= _316;
    end
    always @(posedge _84) begin
        if (_82)
            _322 <= _321;
        else
            _322 <= _319;
    end
    always @(posedge _84) begin
        if (_82)
            _325 <= _324;
        else
            _325 <= _322;
    end
    always @(posedge _84) begin
        if (_82)
            _328 <= _327;
        else
            _328 <= _325;
    end
    assign _357 = _328 & _356;
    assign _358 = _129 & _357;
    assign write_enable_10 = _358 & PHASE_1;
    assign _363 = write_enable_10 | read_enable_8;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_4
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_363), .regcea(vdd), .wea(write_enable_10), .addra(address_10), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_1), .regceb(vdd), .web(write_enable_1), .addrb(address_1), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_370[131:131]), .sbiterrb(_370[130:130]), .doutb(_370[129:66]), .dbiterra(_370[65:65]), .sbiterra(_370[64:64]), .douta(_370[63:0]) );
    assign _371 = _370[63:0];
    assign _301 = ~ PHASE_1;
    assign _7 = _301;
    always @(posedge _84) begin
        if (_82)
            PHASE_1 <= _299;
        else
            if (_72)
                PHASE_1 <= _7;
    end
    assign _383 = PHASE_1 ? _382 : _371;
    assign address_11 = _568 ? _199 : _563;
    assign write_enable_11 = _561 & _568;
    assign address_12 = _568 ? _164 : _68;
    assign _570 = ~ _568;
    assign read_enable_9 = _556 & _570;
    assign _568 = ~ PHASE_4;
    assign write_enable_12 = _554 & _568;
    assign _572 = write_enable_12 | read_enable_9;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_5
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_572), .regcea(vdd), .wea(write_enable_12), .addra(address_12), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_11), .regceb(vdd), .web(write_enable_11), .addrb(address_11), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_577[131:131]), .sbiterrb(_577[130:130]), .doutb(_577[129:66]), .dbiterra(_577[65:65]), .sbiterra(_577[64:64]), .douta(_577[63:0]) );
    assign _578 = _577[63:0];
    assign address_13 = PHASE_4 ? _199 : _563;
    assign _561 = _129 & _524;
    assign write_enable_13 = _561 & PHASE_4;
    assign _486 = _478[129:66];
    assign _485 = _465[129:66];
    assign _487 = PHASE_2 ? _486 : _485;
    assign _483 = _423[129:66];
    assign _482 = _409[129:66];
    assign q1_0 = PHASE_3 ? _483 : _482;
    assign _488 = _390 ? _487 : q1_0;
    assign address_14 = _467 ? _461 : _460;
    assign _473 = ~ _467;
    assign read_enable_10 = _102 & _473;
    assign address_15 = _467 ? _60 : _443;
    assign _469 = ~ _467;
    assign read_enable_11 = _102 & _469;
    assign _467 = ~ PHASE_2;
    assign write_enable_15 = _426 & _467;
    assign _471 = write_enable_15 | read_enable_11;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_6
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_471), .regcea(vdd), .wea(write_enable_15), .addra(address_15), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_10), .regceb(vdd), .web(write_enable_14), .addrb(address_14), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_478[131:131]), .sbiterrb(_478[130:130]), .doutb(_478[129:66]), .dbiterra(_478[65:65]), .sbiterra(_478[64:64]), .douta(_478[63:0]) );
    assign _479 = _478[63:0];
    assign _459 = _172[11:11];
    assign _458 = _172[10:10];
    assign _457 = _172[9:9];
    assign _456 = _172[8:8];
    assign _455 = _172[7:7];
    assign _454 = _172[6:6];
    assign _453 = _172[5:5];
    assign _452 = _172[4:4];
    assign _451 = _172[3:3];
    assign _450 = _172[2:2];
    assign _449 = _172[1:1];
    assign _448 = _172[0:0];
    assign _460 = { _448, _449, _450, _451, _452, _453, _454, _455, _456, _457, _458, _459 };
    assign address_16 = PHASE_2 ? _461 : _460;
    assign _445 = ~ PHASE_2;
    assign read_enable_12 = _102 & _445;
    assign data_13 = wr_d6;
    assign _442 = _137[11:11];
    assign _441 = _137[10:10];
    assign _440 = _137[9:9];
    assign _439 = _137[8:8];
    assign _438 = _137[7:7];
    assign _437 = _137[6:6];
    assign _436 = _137[5:5];
    assign _435 = _137[4:4];
    assign _434 = _137[3:3];
    assign _433 = _137[2:2];
    assign _432 = _137[1:1];
    assign _431 = _137[0:0];
    assign _443 = { _431, _432, _433, _434, _435, _436, _437, _438, _439, _440, _441, _442 };
    assign address_17 = PHASE_2 ? _60 : _443;
    assign _428 = ~ PHASE_2;
    assign read_enable_13 = _102 & _428;
    assign _426 = _62[6:6];
    assign write_enable_17 = _426 & PHASE_2;
    assign _430 = write_enable_17 | read_enable_13;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_7
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_430), .regcea(vdd), .wea(write_enable_17), .addra(address_17), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_12), .regceb(vdd), .web(write_enable_16), .addrb(address_16), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_465[131:131]), .sbiterrb(_465[130:130]), .doutb(_465[129:66]), .dbiterra(_465[65:65]), .sbiterra(_465[64:64]), .douta(_465[63:0]) );
    assign _466 = _465[63:0];
    assign _387 = ~ PHASE_2;
    assign _11 = _387;
    always @(posedge _84) begin
        if (_82)
            PHASE_2 <= _385;
        else
            if (_72)
                PHASE_2 <= _11;
    end
    assign _480 = PHASE_2 ? _479 : _466;
    assign address_18 = _411 ? _199 : _172;
    assign _418 = ~ _411;
    assign read_enable_14 = _102 & _418;
    assign write_enable_18 = _402 & _411;
    assign _420 = write_enable_18 | read_enable_14;
    assign address_19 = _411 ? _164 : _137;
    assign _413 = ~ _411;
    assign read_enable_15 = _102 & _413;
    assign _411 = ~ PHASE_3;
    assign write_enable_19 = _395 & _411;
    assign _415 = write_enable_19 | read_enable_15;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_8
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_415), .regcea(vdd), .wea(write_enable_19), .addra(address_19), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_420), .regceb(vdd), .web(write_enable_18), .addrb(address_18), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_423[131:131]), .sbiterrb(_423[130:130]), .doutb(_423[129:66]), .dbiterra(_423[65:65]), .sbiterra(_423[64:64]), .douta(_423[63:0]) );
    assign _424 = _423[63:0];
    assign _491 = _490[127:64];
    assign data_15 = _491;
    assign address_20 = PHASE_3 ? _199 : _172;
    assign _404 = ~ PHASE_3;
    assign read_enable_16 = _102 & _404;
    assign _401 = ~ _130;
    assign _402 = _129 & _401;
    assign write_enable_20 = _402 & PHASE_3;
    assign _406 = write_enable_20 | read_enable_16;
    assign address_21 = PHASE_3 ? _164 : _137;
    assign _397 = ~ PHASE_3;
    assign read_enable_17 = _102 & _397;
    assign _394 = ~ _130;
    assign _395 = _129 & _394;
    assign write_enable_21 = _395 & PHASE_3;
    assign _399 = write_enable_21 | read_enable_17;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_9
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_399), .regcea(vdd), .wea(write_enable_21), .addra(address_21), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_406), .regceb(vdd), .web(write_enable_20), .addrb(address_20), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_409[131:131]), .sbiterrb(_409[130:130]), .doutb(_409[129:66]), .dbiterra(_409[65:65]), .sbiterra(_409[64:64]), .douta(_409[63:0]) );
    assign _410 = _409[63:0];
    assign _492 = ~ PHASE_3;
    assign _13 = _492;
    always @(posedge _84) begin
        if (_82)
            PHASE_3 <= _392;
        else
            if (_99)
                PHASE_3 <= _13;
    end
    assign q0_0 = PHASE_3 ? _424 : _410;
    always @(posedge _84) begin
        if (_82)
            _390 <= _389;
        else
            _390 <= _92;
    end
    assign _481 = _390 ? _480 : q0_0;
    dp_21
        dp_5
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_481), .d2(_488), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_490[191:128]), .q2(_490[127:64]), .q1(_490[63:0]) );
    assign _493 = _490[63:0];
    assign data_19 = _493;
    assign address_22 = PHASE_4 ? _164 : _68;
    assign _557 = ~ PHASE_4;
    assign _556 = _70[6:6];
    assign read_enable_18 = _556 & _557;
    always @(posedge _84) begin
        if (_82)
            _527 <= _526;
        else
            _527 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _530 <= _529;
        else
            _530 <= _527;
    end
    always @(posedge _84) begin
        if (_82)
            _533 <= _532;
        else
            _533 <= _530;
    end
    always @(posedge _84) begin
        if (_82)
            _536 <= _535;
        else
            _536 <= _533;
    end
    always @(posedge _84) begin
        if (_82)
            _539 <= _538;
        else
            _539 <= _536;
    end
    always @(posedge _84) begin
        if (_82)
            _542 <= _541;
        else
            _542 <= _539;
    end
    always @(posedge _84) begin
        if (_82)
            _545 <= _544;
        else
            _545 <= _542;
    end
    always @(posedge _84) begin
        if (_82)
            _548 <= _547;
        else
            _548 <= _545;
    end
    always @(posedge _84) begin
        if (_82)
            _551 <= _550;
        else
            _551 <= _548;
    end
    assign _552 = ~ _551;
    always @(posedge _84) begin
        if (_82)
            _500 <= _499;
        else
            _500 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _503 <= _502;
        else
            _503 <= _500;
    end
    always @(posedge _84) begin
        if (_82)
            _506 <= _505;
        else
            _506 <= _503;
    end
    always @(posedge _84) begin
        if (_82)
            _509 <= _508;
        else
            _509 <= _506;
    end
    always @(posedge _84) begin
        if (_82)
            _512 <= _511;
        else
            _512 <= _509;
    end
    always @(posedge _84) begin
        if (_82)
            _515 <= _514;
        else
            _515 <= _512;
    end
    always @(posedge _84) begin
        if (_82)
            _518 <= _517;
        else
            _518 <= _515;
    end
    always @(posedge _84) begin
        if (_82)
            _521 <= _520;
        else
            _521 <= _518;
    end
    always @(posedge _84) begin
        if (_82)
            _524 <= _523;
        else
            _524 <= _521;
    end
    assign _553 = _524 & _552;
    assign _554 = _129 & _553;
    assign write_enable_22 = _554 & PHASE_4;
    assign _559 = write_enable_22 | read_enable_18;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_10
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_559), .regcea(vdd), .wea(write_enable_22), .addra(address_22), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_13), .regceb(vdd), .web(write_enable_13), .addrb(address_13), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_566[131:131]), .sbiterrb(_566[130:130]), .doutb(_566[129:66]), .dbiterra(_566[65:65]), .sbiterra(_566[64:64]), .douta(_566[63:0]) );
    assign _567 = _566[63:0];
    assign _497 = ~ PHASE_4;
    assign _15 = _497;
    always @(posedge _84) begin
        if (_82)
            PHASE_4 <= _495;
        else
            if (_72)
                PHASE_4 <= _15;
    end
    assign _579 = PHASE_4 ? _578 : _567;
    assign address_23 = _764 ? _199 : _759;
    assign write_enable_23 = _757 & _764;
    assign address_24 = _764 ? _164 : _68;
    assign _766 = ~ _764;
    assign read_enable_19 = _752 & _766;
    assign _764 = ~ PHASE_7;
    assign write_enable_24 = _750 & _764;
    assign _768 = write_enable_24 | read_enable_19;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_11
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_768), .regcea(vdd), .wea(write_enable_24), .addra(address_24), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_23), .regceb(vdd), .web(write_enable_23), .addrb(address_23), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_773[131:131]), .sbiterrb(_773[130:130]), .doutb(_773[129:66]), .dbiterra(_773[65:65]), .sbiterra(_773[64:64]), .douta(_773[63:0]) );
    assign _774 = _773[63:0];
    assign address_25 = PHASE_7 ? _199 : _759;
    assign _757 = _129 & _720;
    assign write_enable_25 = _757 & PHASE_7;
    assign _682 = _674[129:66];
    assign _681 = _661[129:66];
    assign _683 = PHASE_5 ? _682 : _681;
    assign _679 = _619[129:66];
    assign _678 = _605[129:66];
    assign q1_1 = PHASE_6 ? _679 : _678;
    assign _684 = _586 ? _683 : q1_1;
    assign address_26 = _663 ? _657 : _656;
    assign _669 = ~ _663;
    assign read_enable_20 = _102 & _669;
    assign address_27 = _663 ? _60 : _639;
    assign _665 = ~ _663;
    assign read_enable_21 = _102 & _665;
    assign _663 = ~ PHASE_5;
    assign write_enable_27 = _622 & _663;
    assign _667 = write_enable_27 | read_enable_21;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_12
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_667), .regcea(vdd), .wea(write_enable_27), .addra(address_27), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_20), .regceb(vdd), .web(write_enable_26), .addrb(address_26), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_674[131:131]), .sbiterrb(_674[130:130]), .doutb(_674[129:66]), .dbiterra(_674[65:65]), .sbiterra(_674[64:64]), .douta(_674[63:0]) );
    assign _675 = _674[63:0];
    assign _655 = _172[11:11];
    assign _654 = _172[10:10];
    assign _653 = _172[9:9];
    assign _652 = _172[8:8];
    assign _651 = _172[7:7];
    assign _650 = _172[6:6];
    assign _649 = _172[5:5];
    assign _648 = _172[4:4];
    assign _647 = _172[3:3];
    assign _646 = _172[2:2];
    assign _645 = _172[1:1];
    assign _644 = _172[0:0];
    assign _656 = { _644, _645, _646, _647, _648, _649, _650, _651, _652, _653, _654, _655 };
    assign address_28 = PHASE_5 ? _657 : _656;
    assign _641 = ~ PHASE_5;
    assign read_enable_22 = _102 & _641;
    assign data_25 = wr_d5;
    assign _638 = _137[11:11];
    assign _637 = _137[10:10];
    assign _636 = _137[9:9];
    assign _635 = _137[8:8];
    assign _634 = _137[7:7];
    assign _633 = _137[6:6];
    assign _632 = _137[5:5];
    assign _631 = _137[4:4];
    assign _630 = _137[3:3];
    assign _629 = _137[2:2];
    assign _628 = _137[1:1];
    assign _627 = _137[0:0];
    assign _639 = { _627, _628, _629, _630, _631, _632, _633, _634, _635, _636, _637, _638 };
    assign address_29 = PHASE_5 ? _60 : _639;
    assign _624 = ~ PHASE_5;
    assign read_enable_23 = _102 & _624;
    assign _622 = _62[5:5];
    assign write_enable_29 = _622 & PHASE_5;
    assign _626 = write_enable_29 | read_enable_23;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_13
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_626), .regcea(vdd), .wea(write_enable_29), .addra(address_29), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_22), .regceb(vdd), .web(write_enable_28), .addrb(address_28), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_661[131:131]), .sbiterrb(_661[130:130]), .doutb(_661[129:66]), .dbiterra(_661[65:65]), .sbiterra(_661[64:64]), .douta(_661[63:0]) );
    assign _662 = _661[63:0];
    assign _583 = ~ PHASE_5;
    assign _19 = _583;
    always @(posedge _84) begin
        if (_82)
            PHASE_5 <= _581;
        else
            if (_72)
                PHASE_5 <= _19;
    end
    assign _676 = PHASE_5 ? _675 : _662;
    assign address_30 = _607 ? _199 : _172;
    assign _614 = ~ _607;
    assign read_enable_24 = _102 & _614;
    assign write_enable_30 = _598 & _607;
    assign _616 = write_enable_30 | read_enable_24;
    assign address_31 = _607 ? _164 : _137;
    assign _609 = ~ _607;
    assign read_enable_25 = _102 & _609;
    assign _607 = ~ PHASE_6;
    assign write_enable_31 = _591 & _607;
    assign _611 = write_enable_31 | read_enable_25;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_14
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_611), .regcea(vdd), .wea(write_enable_31), .addra(address_31), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_616), .regceb(vdd), .web(write_enable_30), .addrb(address_30), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_619[131:131]), .sbiterrb(_619[130:130]), .doutb(_619[129:66]), .dbiterra(_619[65:65]), .sbiterra(_619[64:64]), .douta(_619[63:0]) );
    assign _620 = _619[63:0];
    assign _687 = _686[127:64];
    assign data_27 = _687;
    assign address_32 = PHASE_6 ? _199 : _172;
    assign _600 = ~ PHASE_6;
    assign read_enable_26 = _102 & _600;
    assign _597 = ~ _130;
    assign _598 = _129 & _597;
    assign write_enable_32 = _598 & PHASE_6;
    assign _602 = write_enable_32 | read_enable_26;
    assign address_33 = PHASE_6 ? _164 : _137;
    assign _593 = ~ PHASE_6;
    assign read_enable_27 = _102 & _593;
    assign _590 = ~ _130;
    assign _591 = _129 & _590;
    assign write_enable_33 = _591 & PHASE_6;
    assign _595 = write_enable_33 | read_enable_27;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_15
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_595), .regcea(vdd), .wea(write_enable_33), .addra(address_33), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_602), .regceb(vdd), .web(write_enable_32), .addrb(address_32), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_605[131:131]), .sbiterrb(_605[130:130]), .doutb(_605[129:66]), .dbiterra(_605[65:65]), .sbiterra(_605[64:64]), .douta(_605[63:0]) );
    assign _606 = _605[63:0];
    assign _688 = ~ PHASE_6;
    assign _21 = _688;
    always @(posedge _84) begin
        if (_82)
            PHASE_6 <= _588;
        else
            if (_99)
                PHASE_6 <= _21;
    end
    assign q0_1 = PHASE_6 ? _620 : _606;
    always @(posedge _84) begin
        if (_82)
            _586 <= _585;
        else
            _586 <= _92;
    end
    assign _677 = _586 ? _676 : q0_1;
    dp_20
        dp_4
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_677), .d2(_684), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_686[191:128]), .q2(_686[127:64]), .q1(_686[63:0]) );
    assign _689 = _686[63:0];
    assign data_31 = _689;
    assign address_34 = PHASE_7 ? _164 : _68;
    assign _753 = ~ PHASE_7;
    assign _752 = _70[5:5];
    assign read_enable_28 = _752 & _753;
    always @(posedge _84) begin
        if (_82)
            _723 <= _722;
        else
            _723 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _726 <= _725;
        else
            _726 <= _723;
    end
    always @(posedge _84) begin
        if (_82)
            _729 <= _728;
        else
            _729 <= _726;
    end
    always @(posedge _84) begin
        if (_82)
            _732 <= _731;
        else
            _732 <= _729;
    end
    always @(posedge _84) begin
        if (_82)
            _735 <= _734;
        else
            _735 <= _732;
    end
    always @(posedge _84) begin
        if (_82)
            _738 <= _737;
        else
            _738 <= _735;
    end
    always @(posedge _84) begin
        if (_82)
            _741 <= _740;
        else
            _741 <= _738;
    end
    always @(posedge _84) begin
        if (_82)
            _744 <= _743;
        else
            _744 <= _741;
    end
    always @(posedge _84) begin
        if (_82)
            _747 <= _746;
        else
            _747 <= _744;
    end
    assign _748 = ~ _747;
    always @(posedge _84) begin
        if (_82)
            _696 <= _695;
        else
            _696 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _699 <= _698;
        else
            _699 <= _696;
    end
    always @(posedge _84) begin
        if (_82)
            _702 <= _701;
        else
            _702 <= _699;
    end
    always @(posedge _84) begin
        if (_82)
            _705 <= _704;
        else
            _705 <= _702;
    end
    always @(posedge _84) begin
        if (_82)
            _708 <= _707;
        else
            _708 <= _705;
    end
    always @(posedge _84) begin
        if (_82)
            _711 <= _710;
        else
            _711 <= _708;
    end
    always @(posedge _84) begin
        if (_82)
            _714 <= _713;
        else
            _714 <= _711;
    end
    always @(posedge _84) begin
        if (_82)
            _717 <= _716;
        else
            _717 <= _714;
    end
    always @(posedge _84) begin
        if (_82)
            _720 <= _719;
        else
            _720 <= _717;
    end
    assign _749 = _720 & _748;
    assign _750 = _129 & _749;
    assign write_enable_34 = _750 & PHASE_7;
    assign _755 = write_enable_34 | read_enable_28;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_16
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_755), .regcea(vdd), .wea(write_enable_34), .addra(address_34), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_25), .regceb(vdd), .web(write_enable_25), .addrb(address_25), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_762[131:131]), .sbiterrb(_762[130:130]), .doutb(_762[129:66]), .dbiterra(_762[65:65]), .sbiterra(_762[64:64]), .douta(_762[63:0]) );
    assign _763 = _762[63:0];
    assign _693 = ~ PHASE_7;
    assign _23 = _693;
    always @(posedge _84) begin
        if (_82)
            PHASE_7 <= _691;
        else
            if (_72)
                PHASE_7 <= _23;
    end
    assign _775 = PHASE_7 ? _774 : _763;
    assign address_35 = _960 ? _199 : _955;
    assign write_enable_35 = _953 & _960;
    assign address_36 = _960 ? _164 : _68;
    assign _962 = ~ _960;
    assign read_enable_29 = _948 & _962;
    assign _960 = ~ PHASE_10;
    assign write_enable_36 = _946 & _960;
    assign _964 = write_enable_36 | read_enable_29;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_17
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_964), .regcea(vdd), .wea(write_enable_36), .addra(address_36), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_35), .regceb(vdd), .web(write_enable_35), .addrb(address_35), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_969[131:131]), .sbiterrb(_969[130:130]), .doutb(_969[129:66]), .dbiterra(_969[65:65]), .sbiterra(_969[64:64]), .douta(_969[63:0]) );
    assign _970 = _969[63:0];
    assign address_37 = PHASE_10 ? _199 : _955;
    assign _953 = _129 & _916;
    assign write_enable_37 = _953 & PHASE_10;
    assign _878 = _870[129:66];
    assign _877 = _857[129:66];
    assign _879 = PHASE_8 ? _878 : _877;
    assign _875 = _815[129:66];
    assign _874 = _801[129:66];
    assign q1_2 = PHASE_9 ? _875 : _874;
    assign _880 = _782 ? _879 : q1_2;
    assign address_38 = _859 ? _853 : _852;
    assign _865 = ~ _859;
    assign read_enable_30 = _102 & _865;
    assign address_39 = _859 ? _60 : _835;
    assign _861 = ~ _859;
    assign read_enable_31 = _102 & _861;
    assign _859 = ~ PHASE_8;
    assign write_enable_39 = _818 & _859;
    assign _863 = write_enable_39 | read_enable_31;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_18
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_863), .regcea(vdd), .wea(write_enable_39), .addra(address_39), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_30), .regceb(vdd), .web(write_enable_38), .addrb(address_38), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_870[131:131]), .sbiterrb(_870[130:130]), .doutb(_870[129:66]), .dbiterra(_870[65:65]), .sbiterra(_870[64:64]), .douta(_870[63:0]) );
    assign _871 = _870[63:0];
    assign _851 = _172[11:11];
    assign _850 = _172[10:10];
    assign _849 = _172[9:9];
    assign _848 = _172[8:8];
    assign _847 = _172[7:7];
    assign _846 = _172[6:6];
    assign _845 = _172[5:5];
    assign _844 = _172[4:4];
    assign _843 = _172[3:3];
    assign _842 = _172[2:2];
    assign _841 = _172[1:1];
    assign _840 = _172[0:0];
    assign _852 = { _840, _841, _842, _843, _844, _845, _846, _847, _848, _849, _850, _851 };
    assign address_40 = PHASE_8 ? _853 : _852;
    assign _837 = ~ PHASE_8;
    assign read_enable_32 = _102 & _837;
    assign data_37 = wr_d4;
    assign _834 = _137[11:11];
    assign _833 = _137[10:10];
    assign _832 = _137[9:9];
    assign _831 = _137[8:8];
    assign _830 = _137[7:7];
    assign _829 = _137[6:6];
    assign _828 = _137[5:5];
    assign _827 = _137[4:4];
    assign _826 = _137[3:3];
    assign _825 = _137[2:2];
    assign _824 = _137[1:1];
    assign _823 = _137[0:0];
    assign _835 = { _823, _824, _825, _826, _827, _828, _829, _830, _831, _832, _833, _834 };
    assign address_41 = PHASE_8 ? _60 : _835;
    assign _820 = ~ PHASE_8;
    assign read_enable_33 = _102 & _820;
    assign _818 = _62[4:4];
    assign write_enable_41 = _818 & PHASE_8;
    assign _822 = write_enable_41 | read_enable_33;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_19
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_822), .regcea(vdd), .wea(write_enable_41), .addra(address_41), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_32), .regceb(vdd), .web(write_enable_40), .addrb(address_40), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_857[131:131]), .sbiterrb(_857[130:130]), .doutb(_857[129:66]), .dbiterra(_857[65:65]), .sbiterra(_857[64:64]), .douta(_857[63:0]) );
    assign _858 = _857[63:0];
    assign _779 = ~ PHASE_8;
    assign _27 = _779;
    always @(posedge _84) begin
        if (_82)
            PHASE_8 <= _777;
        else
            if (_72)
                PHASE_8 <= _27;
    end
    assign _872 = PHASE_8 ? _871 : _858;
    assign address_42 = _803 ? _199 : _172;
    assign _810 = ~ _803;
    assign read_enable_34 = _102 & _810;
    assign write_enable_42 = _794 & _803;
    assign _812 = write_enable_42 | read_enable_34;
    assign address_43 = _803 ? _164 : _137;
    assign _805 = ~ _803;
    assign read_enable_35 = _102 & _805;
    assign _803 = ~ PHASE_9;
    assign write_enable_43 = _787 & _803;
    assign _807 = write_enable_43 | read_enable_35;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_20
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_807), .regcea(vdd), .wea(write_enable_43), .addra(address_43), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_812), .regceb(vdd), .web(write_enable_42), .addrb(address_42), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_815[131:131]), .sbiterrb(_815[130:130]), .doutb(_815[129:66]), .dbiterra(_815[65:65]), .sbiterra(_815[64:64]), .douta(_815[63:0]) );
    assign _816 = _815[63:0];
    assign _883 = _882[127:64];
    assign data_39 = _883;
    assign address_44 = PHASE_9 ? _199 : _172;
    assign _796 = ~ PHASE_9;
    assign read_enable_36 = _102 & _796;
    assign _793 = ~ _130;
    assign _794 = _129 & _793;
    assign write_enable_44 = _794 & PHASE_9;
    assign _798 = write_enable_44 | read_enable_36;
    assign address_45 = PHASE_9 ? _164 : _137;
    assign _789 = ~ PHASE_9;
    assign read_enable_37 = _102 & _789;
    assign _786 = ~ _130;
    assign _787 = _129 & _786;
    assign write_enable_45 = _787 & PHASE_9;
    assign _791 = write_enable_45 | read_enable_37;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_21
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_791), .regcea(vdd), .wea(write_enable_45), .addra(address_45), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_798), .regceb(vdd), .web(write_enable_44), .addrb(address_44), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_801[131:131]), .sbiterrb(_801[130:130]), .doutb(_801[129:66]), .dbiterra(_801[65:65]), .sbiterra(_801[64:64]), .douta(_801[63:0]) );
    assign _802 = _801[63:0];
    assign _884 = ~ PHASE_9;
    assign _29 = _884;
    always @(posedge _84) begin
        if (_82)
            PHASE_9 <= _784;
        else
            if (_99)
                PHASE_9 <= _29;
    end
    assign q0_2 = PHASE_9 ? _816 : _802;
    always @(posedge _84) begin
        if (_82)
            _782 <= _781;
        else
            _782 <= _92;
    end
    assign _873 = _782 ? _872 : q0_2;
    dp_19
        dp_3
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_873), .d2(_880), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_882[191:128]), .q2(_882[127:64]), .q1(_882[63:0]) );
    assign _885 = _882[63:0];
    assign data_43 = _885;
    assign address_46 = PHASE_10 ? _164 : _68;
    assign _949 = ~ PHASE_10;
    assign _948 = _70[4:4];
    assign read_enable_38 = _948 & _949;
    always @(posedge _84) begin
        if (_82)
            _919 <= _918;
        else
            _919 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _922 <= _921;
        else
            _922 <= _919;
    end
    always @(posedge _84) begin
        if (_82)
            _925 <= _924;
        else
            _925 <= _922;
    end
    always @(posedge _84) begin
        if (_82)
            _928 <= _927;
        else
            _928 <= _925;
    end
    always @(posedge _84) begin
        if (_82)
            _931 <= _930;
        else
            _931 <= _928;
    end
    always @(posedge _84) begin
        if (_82)
            _934 <= _933;
        else
            _934 <= _931;
    end
    always @(posedge _84) begin
        if (_82)
            _937 <= _936;
        else
            _937 <= _934;
    end
    always @(posedge _84) begin
        if (_82)
            _940 <= _939;
        else
            _940 <= _937;
    end
    always @(posedge _84) begin
        if (_82)
            _943 <= _942;
        else
            _943 <= _940;
    end
    assign _944 = ~ _943;
    always @(posedge _84) begin
        if (_82)
            _892 <= _891;
        else
            _892 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _895 <= _894;
        else
            _895 <= _892;
    end
    always @(posedge _84) begin
        if (_82)
            _898 <= _897;
        else
            _898 <= _895;
    end
    always @(posedge _84) begin
        if (_82)
            _901 <= _900;
        else
            _901 <= _898;
    end
    always @(posedge _84) begin
        if (_82)
            _904 <= _903;
        else
            _904 <= _901;
    end
    always @(posedge _84) begin
        if (_82)
            _907 <= _906;
        else
            _907 <= _904;
    end
    always @(posedge _84) begin
        if (_82)
            _910 <= _909;
        else
            _910 <= _907;
    end
    always @(posedge _84) begin
        if (_82)
            _913 <= _912;
        else
            _913 <= _910;
    end
    always @(posedge _84) begin
        if (_82)
            _916 <= _915;
        else
            _916 <= _913;
    end
    assign _945 = _916 & _944;
    assign _946 = _129 & _945;
    assign write_enable_46 = _946 & PHASE_10;
    assign _951 = write_enable_46 | read_enable_38;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_22
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_951), .regcea(vdd), .wea(write_enable_46), .addra(address_46), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_37), .regceb(vdd), .web(write_enable_37), .addrb(address_37), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_958[131:131]), .sbiterrb(_958[130:130]), .doutb(_958[129:66]), .dbiterra(_958[65:65]), .sbiterra(_958[64:64]), .douta(_958[63:0]) );
    assign _959 = _958[63:0];
    assign _889 = ~ PHASE_10;
    assign _31 = _889;
    always @(posedge _84) begin
        if (_82)
            PHASE_10 <= _887;
        else
            if (_72)
                PHASE_10 <= _31;
    end
    assign _971 = PHASE_10 ? _970 : _959;
    assign address_47 = _1156 ? _199 : _1151;
    assign write_enable_47 = _1149 & _1156;
    assign address_48 = _1156 ? _164 : _68;
    assign _1158 = ~ _1156;
    assign read_enable_39 = _1144 & _1158;
    assign _1156 = ~ PHASE_13;
    assign write_enable_48 = _1142 & _1156;
    assign _1160 = write_enable_48 | read_enable_39;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_23
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1160), .regcea(vdd), .wea(write_enable_48), .addra(address_48), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_47), .regceb(vdd), .web(write_enable_47), .addrb(address_47), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1165[131:131]), .sbiterrb(_1165[130:130]), .doutb(_1165[129:66]), .dbiterra(_1165[65:65]), .sbiterra(_1165[64:64]), .douta(_1165[63:0]) );
    assign _1166 = _1165[63:0];
    assign address_49 = PHASE_13 ? _199 : _1151;
    assign _1149 = _129 & _1112;
    assign write_enable_49 = _1149 & PHASE_13;
    assign _1074 = _1066[129:66];
    assign _1073 = _1053[129:66];
    assign _1075 = PHASE_11 ? _1074 : _1073;
    assign _1071 = _1011[129:66];
    assign _1070 = _997[129:66];
    assign q1_3 = PHASE_12 ? _1071 : _1070;
    assign _1076 = _978 ? _1075 : q1_3;
    assign address_50 = _1055 ? _1049 : _1048;
    assign _1061 = ~ _1055;
    assign read_enable_40 = _102 & _1061;
    assign address_51 = _1055 ? _60 : _1031;
    assign _1057 = ~ _1055;
    assign read_enable_41 = _102 & _1057;
    assign _1055 = ~ PHASE_11;
    assign write_enable_51 = _1014 & _1055;
    assign _1059 = write_enable_51 | read_enable_41;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_24
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1059), .regcea(vdd), .wea(write_enable_51), .addra(address_51), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_40), .regceb(vdd), .web(write_enable_50), .addrb(address_50), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1066[131:131]), .sbiterrb(_1066[130:130]), .doutb(_1066[129:66]), .dbiterra(_1066[65:65]), .sbiterra(_1066[64:64]), .douta(_1066[63:0]) );
    assign _1067 = _1066[63:0];
    assign _1047 = _172[11:11];
    assign _1046 = _172[10:10];
    assign _1045 = _172[9:9];
    assign _1044 = _172[8:8];
    assign _1043 = _172[7:7];
    assign _1042 = _172[6:6];
    assign _1041 = _172[5:5];
    assign _1040 = _172[4:4];
    assign _1039 = _172[3:3];
    assign _1038 = _172[2:2];
    assign _1037 = _172[1:1];
    assign _1036 = _172[0:0];
    assign _1048 = { _1036, _1037, _1038, _1039, _1040, _1041, _1042, _1043, _1044, _1045, _1046, _1047 };
    assign address_52 = PHASE_11 ? _1049 : _1048;
    assign _1033 = ~ PHASE_11;
    assign read_enable_42 = _102 & _1033;
    assign data_49 = wr_d3;
    assign _1030 = _137[11:11];
    assign _1029 = _137[10:10];
    assign _1028 = _137[9:9];
    assign _1027 = _137[8:8];
    assign _1026 = _137[7:7];
    assign _1025 = _137[6:6];
    assign _1024 = _137[5:5];
    assign _1023 = _137[4:4];
    assign _1022 = _137[3:3];
    assign _1021 = _137[2:2];
    assign _1020 = _137[1:1];
    assign _1019 = _137[0:0];
    assign _1031 = { _1019, _1020, _1021, _1022, _1023, _1024, _1025, _1026, _1027, _1028, _1029, _1030 };
    assign address_53 = PHASE_11 ? _60 : _1031;
    assign _1016 = ~ PHASE_11;
    assign read_enable_43 = _102 & _1016;
    assign _1014 = _62[3:3];
    assign write_enable_53 = _1014 & PHASE_11;
    assign _1018 = write_enable_53 | read_enable_43;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_25
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1018), .regcea(vdd), .wea(write_enable_53), .addra(address_53), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_42), .regceb(vdd), .web(write_enable_52), .addrb(address_52), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1053[131:131]), .sbiterrb(_1053[130:130]), .doutb(_1053[129:66]), .dbiterra(_1053[65:65]), .sbiterra(_1053[64:64]), .douta(_1053[63:0]) );
    assign _1054 = _1053[63:0];
    assign _975 = ~ PHASE_11;
    assign _35 = _975;
    always @(posedge _84) begin
        if (_82)
            PHASE_11 <= _973;
        else
            if (_72)
                PHASE_11 <= _35;
    end
    assign _1068 = PHASE_11 ? _1067 : _1054;
    assign address_54 = _999 ? _199 : _172;
    assign _1006 = ~ _999;
    assign read_enable_44 = _102 & _1006;
    assign write_enable_54 = _990 & _999;
    assign _1008 = write_enable_54 | read_enable_44;
    assign address_55 = _999 ? _164 : _137;
    assign _1001 = ~ _999;
    assign read_enable_45 = _102 & _1001;
    assign _999 = ~ PHASE_12;
    assign write_enable_55 = _983 & _999;
    assign _1003 = write_enable_55 | read_enable_45;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_26
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1003), .regcea(vdd), .wea(write_enable_55), .addra(address_55), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1008), .regceb(vdd), .web(write_enable_54), .addrb(address_54), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1011[131:131]), .sbiterrb(_1011[130:130]), .doutb(_1011[129:66]), .dbiterra(_1011[65:65]), .sbiterra(_1011[64:64]), .douta(_1011[63:0]) );
    assign _1012 = _1011[63:0];
    assign _1079 = _1078[127:64];
    assign data_51 = _1079;
    assign address_56 = PHASE_12 ? _199 : _172;
    assign _992 = ~ PHASE_12;
    assign read_enable_46 = _102 & _992;
    assign _989 = ~ _130;
    assign _990 = _129 & _989;
    assign write_enable_56 = _990 & PHASE_12;
    assign _994 = write_enable_56 | read_enable_46;
    assign address_57 = PHASE_12 ? _164 : _137;
    assign _985 = ~ PHASE_12;
    assign read_enable_47 = _102 & _985;
    assign _982 = ~ _130;
    assign _983 = _129 & _982;
    assign write_enable_57 = _983 & PHASE_12;
    assign _987 = write_enable_57 | read_enable_47;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_27
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_987), .regcea(vdd), .wea(write_enable_57), .addra(address_57), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_994), .regceb(vdd), .web(write_enable_56), .addrb(address_56), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_997[131:131]), .sbiterrb(_997[130:130]), .doutb(_997[129:66]), .dbiterra(_997[65:65]), .sbiterra(_997[64:64]), .douta(_997[63:0]) );
    assign _998 = _997[63:0];
    assign _1080 = ~ PHASE_12;
    assign _37 = _1080;
    always @(posedge _84) begin
        if (_82)
            PHASE_12 <= _980;
        else
            if (_99)
                PHASE_12 <= _37;
    end
    assign q0_3 = PHASE_12 ? _1012 : _998;
    always @(posedge _84) begin
        if (_82)
            _978 <= _977;
        else
            _978 <= _92;
    end
    assign _1069 = _978 ? _1068 : q0_3;
    dp_18
        dp_2
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1069), .d2(_1076), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1078[191:128]), .q2(_1078[127:64]), .q1(_1078[63:0]) );
    assign _1081 = _1078[63:0];
    assign data_55 = _1081;
    assign address_58 = PHASE_13 ? _164 : _68;
    assign _1145 = ~ PHASE_13;
    assign _1144 = _70[3:3];
    assign read_enable_48 = _1144 & _1145;
    always @(posedge _84) begin
        if (_82)
            _1115 <= _1114;
        else
            _1115 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1118 <= _1117;
        else
            _1118 <= _1115;
    end
    always @(posedge _84) begin
        if (_82)
            _1121 <= _1120;
        else
            _1121 <= _1118;
    end
    always @(posedge _84) begin
        if (_82)
            _1124 <= _1123;
        else
            _1124 <= _1121;
    end
    always @(posedge _84) begin
        if (_82)
            _1127 <= _1126;
        else
            _1127 <= _1124;
    end
    always @(posedge _84) begin
        if (_82)
            _1130 <= _1129;
        else
            _1130 <= _1127;
    end
    always @(posedge _84) begin
        if (_82)
            _1133 <= _1132;
        else
            _1133 <= _1130;
    end
    always @(posedge _84) begin
        if (_82)
            _1136 <= _1135;
        else
            _1136 <= _1133;
    end
    always @(posedge _84) begin
        if (_82)
            _1139 <= _1138;
        else
            _1139 <= _1136;
    end
    assign _1140 = ~ _1139;
    always @(posedge _84) begin
        if (_82)
            _1088 <= _1087;
        else
            _1088 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1091 <= _1090;
        else
            _1091 <= _1088;
    end
    always @(posedge _84) begin
        if (_82)
            _1094 <= _1093;
        else
            _1094 <= _1091;
    end
    always @(posedge _84) begin
        if (_82)
            _1097 <= _1096;
        else
            _1097 <= _1094;
    end
    always @(posedge _84) begin
        if (_82)
            _1100 <= _1099;
        else
            _1100 <= _1097;
    end
    always @(posedge _84) begin
        if (_82)
            _1103 <= _1102;
        else
            _1103 <= _1100;
    end
    always @(posedge _84) begin
        if (_82)
            _1106 <= _1105;
        else
            _1106 <= _1103;
    end
    always @(posedge _84) begin
        if (_82)
            _1109 <= _1108;
        else
            _1109 <= _1106;
    end
    always @(posedge _84) begin
        if (_82)
            _1112 <= _1111;
        else
            _1112 <= _1109;
    end
    assign _1141 = _1112 & _1140;
    assign _1142 = _129 & _1141;
    assign write_enable_58 = _1142 & PHASE_13;
    assign _1147 = write_enable_58 | read_enable_48;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_28
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1147), .regcea(vdd), .wea(write_enable_58), .addra(address_58), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_49), .regceb(vdd), .web(write_enable_49), .addrb(address_49), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1154[131:131]), .sbiterrb(_1154[130:130]), .doutb(_1154[129:66]), .dbiterra(_1154[65:65]), .sbiterra(_1154[64:64]), .douta(_1154[63:0]) );
    assign _1155 = _1154[63:0];
    assign _1085 = ~ PHASE_13;
    assign _39 = _1085;
    always @(posedge _84) begin
        if (_82)
            PHASE_13 <= _1083;
        else
            if (_72)
                PHASE_13 <= _39;
    end
    assign _1167 = PHASE_13 ? _1166 : _1155;
    assign address_59 = _1352 ? _199 : _1347;
    assign write_enable_59 = _1345 & _1352;
    assign address_60 = _1352 ? _164 : _68;
    assign _1354 = ~ _1352;
    assign read_enable_49 = _1340 & _1354;
    assign _1352 = ~ PHASE_16;
    assign write_enable_60 = _1338 & _1352;
    assign _1356 = write_enable_60 | read_enable_49;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_29
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1356), .regcea(vdd), .wea(write_enable_60), .addra(address_60), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_59), .regceb(vdd), .web(write_enable_59), .addrb(address_59), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1361[131:131]), .sbiterrb(_1361[130:130]), .doutb(_1361[129:66]), .dbiterra(_1361[65:65]), .sbiterra(_1361[64:64]), .douta(_1361[63:0]) );
    assign _1362 = _1361[63:0];
    assign address_61 = PHASE_16 ? _199 : _1347;
    assign _1345 = _129 & _1308;
    assign write_enable_61 = _1345 & PHASE_16;
    assign _1270 = _1262[129:66];
    assign _1269 = _1249[129:66];
    assign _1271 = PHASE_14 ? _1270 : _1269;
    assign _1267 = _1207[129:66];
    assign _1266 = _1193[129:66];
    assign q1_4 = PHASE_15 ? _1267 : _1266;
    assign _1272 = _1174 ? _1271 : q1_4;
    assign address_62 = _1251 ? _1245 : _1244;
    assign _1257 = ~ _1251;
    assign read_enable_50 = _102 & _1257;
    assign address_63 = _1251 ? _60 : _1227;
    assign _1253 = ~ _1251;
    assign read_enable_51 = _102 & _1253;
    assign _1251 = ~ PHASE_14;
    assign write_enable_63 = _1210 & _1251;
    assign _1255 = write_enable_63 | read_enable_51;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_30
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1255), .regcea(vdd), .wea(write_enable_63), .addra(address_63), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_50), .regceb(vdd), .web(write_enable_62), .addrb(address_62), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1262[131:131]), .sbiterrb(_1262[130:130]), .doutb(_1262[129:66]), .dbiterra(_1262[65:65]), .sbiterra(_1262[64:64]), .douta(_1262[63:0]) );
    assign _1263 = _1262[63:0];
    assign _1243 = _172[11:11];
    assign _1242 = _172[10:10];
    assign _1241 = _172[9:9];
    assign _1240 = _172[8:8];
    assign _1239 = _172[7:7];
    assign _1238 = _172[6:6];
    assign _1237 = _172[5:5];
    assign _1236 = _172[4:4];
    assign _1235 = _172[3:3];
    assign _1234 = _172[2:2];
    assign _1233 = _172[1:1];
    assign _1232 = _172[0:0];
    assign _1244 = { _1232, _1233, _1234, _1235, _1236, _1237, _1238, _1239, _1240, _1241, _1242, _1243 };
    assign address_64 = PHASE_14 ? _1245 : _1244;
    assign _1229 = ~ PHASE_14;
    assign read_enable_52 = _102 & _1229;
    assign data_61 = wr_d2;
    assign _1226 = _137[11:11];
    assign _1225 = _137[10:10];
    assign _1224 = _137[9:9];
    assign _1223 = _137[8:8];
    assign _1222 = _137[7:7];
    assign _1221 = _137[6:6];
    assign _1220 = _137[5:5];
    assign _1219 = _137[4:4];
    assign _1218 = _137[3:3];
    assign _1217 = _137[2:2];
    assign _1216 = _137[1:1];
    assign _1215 = _137[0:0];
    assign _1227 = { _1215, _1216, _1217, _1218, _1219, _1220, _1221, _1222, _1223, _1224, _1225, _1226 };
    assign address_65 = PHASE_14 ? _60 : _1227;
    assign _1212 = ~ PHASE_14;
    assign read_enable_53 = _102 & _1212;
    assign _1210 = _62[2:2];
    assign write_enable_65 = _1210 & PHASE_14;
    assign _1214 = write_enable_65 | read_enable_53;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_31
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1214), .regcea(vdd), .wea(write_enable_65), .addra(address_65), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_52), .regceb(vdd), .web(write_enable_64), .addrb(address_64), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1249[131:131]), .sbiterrb(_1249[130:130]), .doutb(_1249[129:66]), .dbiterra(_1249[65:65]), .sbiterra(_1249[64:64]), .douta(_1249[63:0]) );
    assign _1250 = _1249[63:0];
    assign _1171 = ~ PHASE_14;
    assign _43 = _1171;
    always @(posedge _84) begin
        if (_82)
            PHASE_14 <= _1169;
        else
            if (_72)
                PHASE_14 <= _43;
    end
    assign _1264 = PHASE_14 ? _1263 : _1250;
    assign address_66 = _1195 ? _199 : _172;
    assign _1202 = ~ _1195;
    assign read_enable_54 = _102 & _1202;
    assign write_enable_66 = _1186 & _1195;
    assign _1204 = write_enable_66 | read_enable_54;
    assign address_67 = _1195 ? _164 : _137;
    assign _1197 = ~ _1195;
    assign read_enable_55 = _102 & _1197;
    assign _1195 = ~ PHASE_15;
    assign write_enable_67 = _1179 & _1195;
    assign _1199 = write_enable_67 | read_enable_55;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_32
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1199), .regcea(vdd), .wea(write_enable_67), .addra(address_67), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1204), .regceb(vdd), .web(write_enable_66), .addrb(address_66), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1207[131:131]), .sbiterrb(_1207[130:130]), .doutb(_1207[129:66]), .dbiterra(_1207[65:65]), .sbiterra(_1207[64:64]), .douta(_1207[63:0]) );
    assign _1208 = _1207[63:0];
    assign _1275 = _1274[127:64];
    assign data_63 = _1275;
    assign address_68 = PHASE_15 ? _199 : _172;
    assign _1188 = ~ PHASE_15;
    assign read_enable_56 = _102 & _1188;
    assign _1185 = ~ _130;
    assign _1186 = _129 & _1185;
    assign write_enable_68 = _1186 & PHASE_15;
    assign _1190 = write_enable_68 | read_enable_56;
    assign address_69 = PHASE_15 ? _164 : _137;
    assign _1181 = ~ PHASE_15;
    assign read_enable_57 = _102 & _1181;
    assign _1178 = ~ _130;
    assign _1179 = _129 & _1178;
    assign write_enable_69 = _1179 & PHASE_15;
    assign _1183 = write_enable_69 | read_enable_57;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_33
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1183), .regcea(vdd), .wea(write_enable_69), .addra(address_69), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1190), .regceb(vdd), .web(write_enable_68), .addrb(address_68), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1193[131:131]), .sbiterrb(_1193[130:130]), .doutb(_1193[129:66]), .dbiterra(_1193[65:65]), .sbiterra(_1193[64:64]), .douta(_1193[63:0]) );
    assign _1194 = _1193[63:0];
    assign _1276 = ~ PHASE_15;
    assign _45 = _1276;
    always @(posedge _84) begin
        if (_82)
            PHASE_15 <= _1176;
        else
            if (_99)
                PHASE_15 <= _45;
    end
    assign q0_4 = PHASE_15 ? _1208 : _1194;
    always @(posedge _84) begin
        if (_82)
            _1174 <= _1173;
        else
            _1174 <= _92;
    end
    assign _1265 = _1174 ? _1264 : q0_4;
    dp_17
        dp_1
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1265), .d2(_1272), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1274[191:128]), .q2(_1274[127:64]), .q1(_1274[63:0]) );
    assign _1277 = _1274[63:0];
    assign data_67 = _1277;
    assign address_70 = PHASE_16 ? _164 : _68;
    assign _1341 = ~ PHASE_16;
    assign _1340 = _70[2:2];
    assign read_enable_58 = _1340 & _1341;
    always @(posedge _84) begin
        if (_82)
            _1311 <= _1310;
        else
            _1311 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1314 <= _1313;
        else
            _1314 <= _1311;
    end
    always @(posedge _84) begin
        if (_82)
            _1317 <= _1316;
        else
            _1317 <= _1314;
    end
    always @(posedge _84) begin
        if (_82)
            _1320 <= _1319;
        else
            _1320 <= _1317;
    end
    always @(posedge _84) begin
        if (_82)
            _1323 <= _1322;
        else
            _1323 <= _1320;
    end
    always @(posedge _84) begin
        if (_82)
            _1326 <= _1325;
        else
            _1326 <= _1323;
    end
    always @(posedge _84) begin
        if (_82)
            _1329 <= _1328;
        else
            _1329 <= _1326;
    end
    always @(posedge _84) begin
        if (_82)
            _1332 <= _1331;
        else
            _1332 <= _1329;
    end
    always @(posedge _84) begin
        if (_82)
            _1335 <= _1334;
        else
            _1335 <= _1332;
    end
    assign _1336 = ~ _1335;
    always @(posedge _84) begin
        if (_82)
            _1284 <= _1283;
        else
            _1284 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1287 <= _1286;
        else
            _1287 <= _1284;
    end
    always @(posedge _84) begin
        if (_82)
            _1290 <= _1289;
        else
            _1290 <= _1287;
    end
    always @(posedge _84) begin
        if (_82)
            _1293 <= _1292;
        else
            _1293 <= _1290;
    end
    always @(posedge _84) begin
        if (_82)
            _1296 <= _1295;
        else
            _1296 <= _1293;
    end
    always @(posedge _84) begin
        if (_82)
            _1299 <= _1298;
        else
            _1299 <= _1296;
    end
    always @(posedge _84) begin
        if (_82)
            _1302 <= _1301;
        else
            _1302 <= _1299;
    end
    always @(posedge _84) begin
        if (_82)
            _1305 <= _1304;
        else
            _1305 <= _1302;
    end
    always @(posedge _84) begin
        if (_82)
            _1308 <= _1307;
        else
            _1308 <= _1305;
    end
    assign _1337 = _1308 & _1336;
    assign _1338 = _129 & _1337;
    assign write_enable_70 = _1338 & PHASE_16;
    assign _1343 = write_enable_70 | read_enable_58;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_34
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1343), .regcea(vdd), .wea(write_enable_70), .addra(address_70), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_61), .regceb(vdd), .web(write_enable_61), .addrb(address_61), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1350[131:131]), .sbiterrb(_1350[130:130]), .doutb(_1350[129:66]), .dbiterra(_1350[65:65]), .sbiterra(_1350[64:64]), .douta(_1350[63:0]) );
    assign _1351 = _1350[63:0];
    assign _1281 = ~ PHASE_16;
    assign _47 = _1281;
    always @(posedge _84) begin
        if (_82)
            PHASE_16 <= _1279;
        else
            if (_72)
                PHASE_16 <= _47;
    end
    assign _1363 = PHASE_16 ? _1362 : _1351;
    assign address_71 = _1548 ? _199 : _1543;
    assign write_enable_71 = _1541 & _1548;
    assign address_72 = _1548 ? _164 : _68;
    assign _1550 = ~ _1548;
    assign read_enable_59 = _1536 & _1550;
    assign _1548 = ~ PHASE_19;
    assign write_enable_72 = _1534 & _1548;
    assign _1552 = write_enable_72 | read_enable_59;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_35
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1552), .regcea(vdd), .wea(write_enable_72), .addra(address_72), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_71), .regceb(vdd), .web(write_enable_71), .addrb(address_71), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1557[131:131]), .sbiterrb(_1557[130:130]), .doutb(_1557[129:66]), .dbiterra(_1557[65:65]), .sbiterra(_1557[64:64]), .douta(_1557[63:0]) );
    assign _1558 = _1557[63:0];
    assign address_73 = PHASE_19 ? _199 : _1543;
    assign _1541 = _129 & _1504;
    assign write_enable_73 = _1541 & PHASE_19;
    assign _1466 = _1458[129:66];
    assign _1465 = _1445[129:66];
    assign _1467 = PHASE_17 ? _1466 : _1465;
    assign _1463 = _1403[129:66];
    assign _1462 = _1389[129:66];
    assign q1_5 = PHASE_18 ? _1463 : _1462;
    assign _1468 = _1370 ? _1467 : q1_5;
    assign address_74 = _1447 ? _1441 : _1440;
    assign _1453 = ~ _1447;
    assign read_enable_60 = _102 & _1453;
    assign address_75 = _1447 ? _60 : _1423;
    assign _1449 = ~ _1447;
    assign read_enable_61 = _102 & _1449;
    assign _1447 = ~ PHASE_17;
    assign write_enable_75 = _1406 & _1447;
    assign _1451 = write_enable_75 | read_enable_61;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_36
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1451), .regcea(vdd), .wea(write_enable_75), .addra(address_75), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_60), .regceb(vdd), .web(write_enable_74), .addrb(address_74), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1458[131:131]), .sbiterrb(_1458[130:130]), .doutb(_1458[129:66]), .dbiterra(_1458[65:65]), .sbiterra(_1458[64:64]), .douta(_1458[63:0]) );
    assign _1459 = _1458[63:0];
    assign _1439 = _172[11:11];
    assign _1438 = _172[10:10];
    assign _1437 = _172[9:9];
    assign _1436 = _172[8:8];
    assign _1435 = _172[7:7];
    assign _1434 = _172[6:6];
    assign _1433 = _172[5:5];
    assign _1432 = _172[4:4];
    assign _1431 = _172[3:3];
    assign _1430 = _172[2:2];
    assign _1429 = _172[1:1];
    assign _1428 = _172[0:0];
    assign _1440 = { _1428, _1429, _1430, _1431, _1432, _1433, _1434, _1435, _1436, _1437, _1438, _1439 };
    assign address_76 = PHASE_17 ? _1441 : _1440;
    assign _1425 = ~ PHASE_17;
    assign read_enable_62 = _102 & _1425;
    assign data_73 = wr_d1;
    assign _1422 = _137[11:11];
    assign _1421 = _137[10:10];
    assign _1420 = _137[9:9];
    assign _1419 = _137[8:8];
    assign _1418 = _137[7:7];
    assign _1417 = _137[6:6];
    assign _1416 = _137[5:5];
    assign _1415 = _137[4:4];
    assign _1414 = _137[3:3];
    assign _1413 = _137[2:2];
    assign _1412 = _137[1:1];
    assign _1411 = _137[0:0];
    assign _1423 = { _1411, _1412, _1413, _1414, _1415, _1416, _1417, _1418, _1419, _1420, _1421, _1422 };
    assign address_77 = PHASE_17 ? _60 : _1423;
    assign _1408 = ~ PHASE_17;
    assign read_enable_63 = _102 & _1408;
    assign _1406 = _62[1:1];
    assign write_enable_77 = _1406 & PHASE_17;
    assign _1410 = write_enable_77 | read_enable_63;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_37
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1410), .regcea(vdd), .wea(write_enable_77), .addra(address_77), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_62), .regceb(vdd), .web(write_enable_76), .addrb(address_76), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1445[131:131]), .sbiterrb(_1445[130:130]), .doutb(_1445[129:66]), .dbiterra(_1445[65:65]), .sbiterra(_1445[64:64]), .douta(_1445[63:0]) );
    assign _1446 = _1445[63:0];
    assign _1367 = ~ PHASE_17;
    assign _51 = _1367;
    always @(posedge _84) begin
        if (_82)
            PHASE_17 <= _1365;
        else
            if (_72)
                PHASE_17 <= _51;
    end
    assign _1460 = PHASE_17 ? _1459 : _1446;
    assign address_78 = _1391 ? _199 : _172;
    assign _1398 = ~ _1391;
    assign read_enable_64 = _102 & _1398;
    assign write_enable_78 = _1382 & _1391;
    assign _1400 = write_enable_78 | read_enable_64;
    assign address_79 = _1391 ? _164 : _137;
    assign _1393 = ~ _1391;
    assign read_enable_65 = _102 & _1393;
    assign _1391 = ~ PHASE_18;
    assign write_enable_79 = _1375 & _1391;
    assign _1395 = write_enable_79 | read_enable_65;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_38
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1395), .regcea(vdd), .wea(write_enable_79), .addra(address_79), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1400), .regceb(vdd), .web(write_enable_78), .addrb(address_78), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1403[131:131]), .sbiterrb(_1403[130:130]), .doutb(_1403[129:66]), .dbiterra(_1403[65:65]), .sbiterra(_1403[64:64]), .douta(_1403[63:0]) );
    assign _1404 = _1403[63:0];
    assign _1471 = _1470[127:64];
    assign data_75 = _1471;
    assign address_80 = PHASE_18 ? _199 : _172;
    assign _1384 = ~ PHASE_18;
    assign read_enable_66 = _102 & _1384;
    assign _1381 = ~ _130;
    assign _1382 = _129 & _1381;
    assign write_enable_80 = _1382 & PHASE_18;
    assign _1386 = write_enable_80 | read_enable_66;
    assign address_81 = PHASE_18 ? _164 : _137;
    assign _1377 = ~ PHASE_18;
    assign read_enable_67 = _102 & _1377;
    assign _1374 = ~ _130;
    assign _1375 = _129 & _1374;
    assign write_enable_81 = _1375 & PHASE_18;
    assign _1379 = write_enable_81 | read_enable_67;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_39
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1379), .regcea(vdd), .wea(write_enable_81), .addra(address_81), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1386), .regceb(vdd), .web(write_enable_80), .addrb(address_80), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1389[131:131]), .sbiterrb(_1389[130:130]), .doutb(_1389[129:66]), .dbiterra(_1389[65:65]), .sbiterra(_1389[64:64]), .douta(_1389[63:0]) );
    assign _1390 = _1389[63:0];
    assign _1472 = ~ PHASE_18;
    assign _53 = _1472;
    always @(posedge _84) begin
        if (_82)
            PHASE_18 <= _1372;
        else
            if (_99)
                PHASE_18 <= _53;
    end
    assign q0_5 = PHASE_18 ? _1404 : _1390;
    always @(posedge _84) begin
        if (_82)
            _1370 <= _1369;
        else
            _1370 <= _92;
    end
    assign _1461 = _1370 ? _1460 : q0_5;
    dp_16
        dp_0
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1461), .d2(_1468), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1470[191:128]), .q2(_1470[127:64]), .q1(_1470[63:0]) );
    assign _1473 = _1470[63:0];
    assign data_79 = _1473;
    assign address_82 = PHASE_19 ? _164 : _68;
    assign _1537 = ~ PHASE_19;
    assign _1536 = _70[1:1];
    assign read_enable_68 = _1536 & _1537;
    always @(posedge _84) begin
        if (_82)
            _1507 <= _1506;
        else
            _1507 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1510 <= _1509;
        else
            _1510 <= _1507;
    end
    always @(posedge _84) begin
        if (_82)
            _1513 <= _1512;
        else
            _1513 <= _1510;
    end
    always @(posedge _84) begin
        if (_82)
            _1516 <= _1515;
        else
            _1516 <= _1513;
    end
    always @(posedge _84) begin
        if (_82)
            _1519 <= _1518;
        else
            _1519 <= _1516;
    end
    always @(posedge _84) begin
        if (_82)
            _1522 <= _1521;
        else
            _1522 <= _1519;
    end
    always @(posedge _84) begin
        if (_82)
            _1525 <= _1524;
        else
            _1525 <= _1522;
    end
    always @(posedge _84) begin
        if (_82)
            _1528 <= _1527;
        else
            _1528 <= _1525;
    end
    always @(posedge _84) begin
        if (_82)
            _1531 <= _1530;
        else
            _1531 <= _1528;
    end
    assign _1532 = ~ _1531;
    always @(posedge _84) begin
        if (_82)
            _1480 <= _1479;
        else
            _1480 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1483 <= _1482;
        else
            _1483 <= _1480;
    end
    always @(posedge _84) begin
        if (_82)
            _1486 <= _1485;
        else
            _1486 <= _1483;
    end
    always @(posedge _84) begin
        if (_82)
            _1489 <= _1488;
        else
            _1489 <= _1486;
    end
    always @(posedge _84) begin
        if (_82)
            _1492 <= _1491;
        else
            _1492 <= _1489;
    end
    always @(posedge _84) begin
        if (_82)
            _1495 <= _1494;
        else
            _1495 <= _1492;
    end
    always @(posedge _84) begin
        if (_82)
            _1498 <= _1497;
        else
            _1498 <= _1495;
    end
    always @(posedge _84) begin
        if (_82)
            _1501 <= _1500;
        else
            _1501 <= _1498;
    end
    always @(posedge _84) begin
        if (_82)
            _1504 <= _1503;
        else
            _1504 <= _1501;
    end
    assign _1533 = _1504 & _1532;
    assign _1534 = _129 & _1533;
    assign write_enable_82 = _1534 & PHASE_19;
    assign _1539 = write_enable_82 | read_enable_68;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_40
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1539), .regcea(vdd), .wea(write_enable_82), .addra(address_82), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_73), .regceb(vdd), .web(write_enable_73), .addrb(address_73), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1546[131:131]), .sbiterrb(_1546[130:130]), .doutb(_1546[129:66]), .dbiterra(_1546[65:65]), .sbiterra(_1546[64:64]), .douta(_1546[63:0]) );
    assign _1547 = _1546[63:0];
    assign _1477 = ~ PHASE_19;
    assign _55 = _1477;
    always @(posedge _84) begin
        if (_82)
            PHASE_19 <= _1475;
        else
            if (_72)
                PHASE_19 <= _55;
    end
    assign _1559 = PHASE_19 ? _1558 : _1547;
    assign address_83 = _1744 ? _199 : _1739;
    assign write_enable_83 = _1737 & _1744;
    assign address_84 = _1744 ? _164 : _68;
    assign _1746 = ~ _1744;
    assign read_enable_69 = _1732 & _1746;
    assign _1744 = ~ PHASE_22;
    assign write_enable_84 = _1730 & _1744;
    assign _1748 = write_enable_84 | read_enable_69;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_41
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1748), .regcea(vdd), .wea(write_enable_84), .addra(address_84), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_83), .regceb(vdd), .web(write_enable_83), .addrb(address_83), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1753[131:131]), .sbiterrb(_1753[130:130]), .doutb(_1753[129:66]), .dbiterra(_1753[65:65]), .sbiterra(_1753[64:64]), .douta(_1753[63:0]) );
    assign _1754 = _1753[63:0];
    assign address_85 = PHASE_22 ? _199 : _1739;
    assign _1737 = _129 & _1700;
    assign write_enable_85 = _1737 & PHASE_22;
    assign _292 = _91[521:518];
    assign _291 = _91[517:517];
    assign _289 = _91[513:513];
    assign _288 = _91[512:449];
    assign _287 = _91[448:385];
    assign _286 = _91[384:321];
    assign _285 = _91[320:257];
    assign _284 = _91[256:193];
    assign _283 = _91[192:129];
    assign _282 = _91[128:65];
    assign _1662 = _1654[129:66];
    assign _1661 = _1641[129:66];
    assign _1663 = PHASE_20 ? _1662 : _1661;
    assign _1659 = _1599[129:66];
    assign _1658 = _1585[129:66];
    assign q1_6 = PHASE_21 ? _1659 : _1658;
    assign _1664 = _1566 ? _1663 : q1_6;
    assign address_86 = _1643 ? _1637 : _1636;
    assign _1649 = ~ _1643;
    assign read_enable_70 = _102 & _1649;
    assign address_87 = _1643 ? _60 : _1619;
    assign _1645 = ~ _1643;
    assign read_enable_71 = _102 & _1645;
    assign _1643 = ~ PHASE_20;
    assign write_enable_87 = _1602 & _1643;
    assign _1647 = write_enable_87 | read_enable_71;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_42
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1647), .regcea(vdd), .wea(write_enable_87), .addra(address_87), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_70), .regceb(vdd), .web(write_enable_86), .addrb(address_86), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1654[131:131]), .sbiterrb(_1654[130:130]), .doutb(_1654[129:66]), .dbiterra(_1654[65:65]), .sbiterra(_1654[64:64]), .douta(_1654[63:0]) );
    assign _1655 = _1654[63:0];
    assign _1635 = _172[11:11];
    assign _1634 = _172[10:10];
    assign _1633 = _172[9:9];
    assign _1632 = _172[8:8];
    assign _1631 = _172[7:7];
    assign _1630 = _172[6:6];
    assign _1629 = _172[5:5];
    assign _1628 = _172[4:4];
    assign _1627 = _172[3:3];
    assign _1626 = _172[2:2];
    assign _1625 = _172[1:1];
    assign _1624 = _172[0:0];
    assign _1636 = { _1624, _1625, _1626, _1627, _1628, _1629, _1630, _1631, _1632, _1633, _1634, _1635 };
    assign address_88 = PHASE_20 ? _1637 : _1636;
    assign _1621 = ~ PHASE_20;
    assign read_enable_72 = _102 & _1621;
    assign data_85 = wr_d0;
    assign _60 = wr_addr;
    assign _1618 = _137[11:11];
    assign _1617 = _137[10:10];
    assign _1616 = _137[9:9];
    assign _1615 = _137[8:8];
    assign _1614 = _137[7:7];
    assign _1613 = _137[6:6];
    assign _1612 = _137[5:5];
    assign _1611 = _137[4:4];
    assign _1610 = _137[3:3];
    assign _1609 = _137[2:2];
    assign _1608 = _137[1:1];
    assign _1607 = _137[0:0];
    assign _1619 = { _1607, _1608, _1609, _1610, _1611, _1612, _1613, _1614, _1615, _1616, _1617, _1618 };
    assign address_89 = PHASE_20 ? _60 : _1619;
    assign _1604 = ~ PHASE_20;
    assign read_enable_73 = _102 & _1604;
    assign _62 = wr_en;
    assign _1602 = _62[0:0];
    assign write_enable_89 = _1602 & PHASE_20;
    assign _1606 = write_enable_89 | read_enable_73;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_43
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1606), .regcea(vdd), .wea(write_enable_89), .addra(address_89), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_72), .regceb(vdd), .web(write_enable_88), .addrb(address_88), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1641[131:131]), .sbiterrb(_1641[130:130]), .doutb(_1641[129:66]), .dbiterra(_1641[65:65]), .sbiterra(_1641[64:64]), .douta(_1641[63:0]) );
    assign _1642 = _1641[63:0];
    assign _1563 = ~ PHASE_20;
    assign _63 = _1563;
    always @(posedge _84) begin
        if (_82)
            PHASE_20 <= _1561;
        else
            if (_72)
                PHASE_20 <= _63;
    end
    assign _1656 = PHASE_20 ? _1655 : _1642;
    assign address_90 = _1587 ? _199 : _172;
    assign _1594 = ~ _1587;
    assign read_enable_74 = _102 & _1594;
    assign write_enable_90 = _1578 & _1587;
    assign _1596 = write_enable_90 | read_enable_74;
    assign address_91 = _1587 ? _164 : _137;
    assign _1589 = ~ _1587;
    assign read_enable_75 = _102 & _1589;
    assign _1587 = ~ PHASE_21;
    assign write_enable_91 = _1571 & _1587;
    assign _1591 = write_enable_91 | read_enable_75;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_44
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1591), .regcea(vdd), .wea(write_enable_91), .addra(address_91), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1596), .regceb(vdd), .web(write_enable_90), .addrb(address_90), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1599[131:131]), .sbiterrb(_1599[130:130]), .doutb(_1599[129:66]), .dbiterra(_1599[65:65]), .sbiterra(_1599[64:64]), .douta(_1599[63:0]) );
    assign _1600 = _1599[63:0];
    assign _1667 = _1666[127:64];
    assign data_87 = _1667;
    always @(posedge _84) begin
        if (_82)
            _175 <= _174;
        else
            _175 <= _172;
    end
    always @(posedge _84) begin
        if (_82)
            _178 <= _177;
        else
            _178 <= _175;
    end
    always @(posedge _84) begin
        if (_82)
            _181 <= _180;
        else
            _181 <= _178;
    end
    always @(posedge _84) begin
        if (_82)
            _184 <= _183;
        else
            _184 <= _181;
    end
    always @(posedge _84) begin
        if (_82)
            _187 <= _186;
        else
            _187 <= _184;
    end
    always @(posedge _84) begin
        if (_82)
            _190 <= _189;
        else
            _190 <= _187;
    end
    always @(posedge _84) begin
        if (_82)
            _193 <= _192;
        else
            _193 <= _190;
    end
    always @(posedge _84) begin
        if (_82)
            _196 <= _195;
        else
            _196 <= _193;
    end
    always @(posedge _84) begin
        if (_82)
            _199 <= _198;
        else
            _199 <= _196;
    end
    assign _172 = _91[64:53];
    assign address_92 = PHASE_21 ? _199 : _172;
    assign _1580 = ~ PHASE_21;
    assign read_enable_76 = _102 & _1580;
    assign _1577 = ~ _130;
    assign _1578 = _129 & _1577;
    assign write_enable_92 = _1578 & PHASE_21;
    assign _1582 = write_enable_92 | read_enable_76;
    assign address_93 = PHASE_21 ? _164 : _137;
    assign _1573 = ~ PHASE_21;
    assign read_enable_77 = _102 & _1573;
    assign _1570 = ~ _130;
    assign _1571 = _129 & _1570;
    assign write_enable_93 = _1571 & PHASE_21;
    assign _1575 = write_enable_93 | read_enable_77;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_45
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1575), .regcea(vdd), .wea(write_enable_93), .addra(address_93), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1582), .regceb(vdd), .web(write_enable_92), .addrb(address_92), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1585[131:131]), .sbiterrb(_1585[130:130]), .doutb(_1585[129:66]), .dbiterra(_1585[65:65]), .sbiterra(_1585[64:64]), .douta(_1585[63:0]) );
    assign _1586 = _1585[63:0];
    assign _99 = _91[523:523];
    assign _1668 = ~ PHASE_21;
    assign _65 = _1668;
    always @(posedge _84) begin
        if (_82)
            PHASE_21 <= _1568;
        else
            if (_99)
                PHASE_21 <= _65;
    end
    assign q0_6 = PHASE_21 ? _1600 : _1586;
    assign _92 = _91[514:514];
    always @(posedge _84) begin
        if (_82)
            _1566 <= _1565;
        else
            _1566 <= _92;
    end
    assign _1657 = _1566 ? _1656 : q0_6;
    dp_15
        dp
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1657), .d2(_1664), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1666[191:128]), .q2(_1666[127:64]), .q1(_1666[63:0]) );
    assign _1669 = _1666[63:0];
    assign data_91 = _1669;
    assign _137 = _91[52:41];
    always @(posedge _84) begin
        if (_82)
            _140 <= _139;
        else
            _140 <= _137;
    end
    always @(posedge _84) begin
        if (_82)
            _143 <= _142;
        else
            _143 <= _140;
    end
    always @(posedge _84) begin
        if (_82)
            _146 <= _145;
        else
            _146 <= _143;
    end
    always @(posedge _84) begin
        if (_82)
            _149 <= _148;
        else
            _149 <= _146;
    end
    always @(posedge _84) begin
        if (_82)
            _152 <= _151;
        else
            _152 <= _149;
    end
    always @(posedge _84) begin
        if (_82)
            _155 <= _154;
        else
            _155 <= _152;
    end
    always @(posedge _84) begin
        if (_82)
            _158 <= _157;
        else
            _158 <= _155;
    end
    always @(posedge _84) begin
        if (_82)
            _161 <= _160;
        else
            _161 <= _158;
    end
    always @(posedge _84) begin
        if (_82)
            _164 <= _163;
        else
            _164 <= _161;
    end
    assign _68 = rd_addr;
    assign address_94 = PHASE_22 ? _164 : _68;
    assign _1733 = ~ PHASE_22;
    assign _70 = rd_en;
    assign _1732 = _70[0:0];
    assign read_enable_78 = _1732 & _1733;
    assign _290 = _91[516:516];
    always @(posedge _84) begin
        if (_82)
            _1703 <= _1702;
        else
            _1703 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1706 <= _1705;
        else
            _1706 <= _1703;
    end
    always @(posedge _84) begin
        if (_82)
            _1709 <= _1708;
        else
            _1709 <= _1706;
    end
    always @(posedge _84) begin
        if (_82)
            _1712 <= _1711;
        else
            _1712 <= _1709;
    end
    always @(posedge _84) begin
        if (_82)
            _1715 <= _1714;
        else
            _1715 <= _1712;
    end
    always @(posedge _84) begin
        if (_82)
            _1718 <= _1717;
        else
            _1718 <= _1715;
    end
    always @(posedge _84) begin
        if (_82)
            _1721 <= _1720;
        else
            _1721 <= _1718;
    end
    always @(posedge _84) begin
        if (_82)
            _1724 <= _1723;
        else
            _1724 <= _1721;
    end
    always @(posedge _84) begin
        if (_82)
            _1727 <= _1726;
        else
            _1727 <= _1724;
    end
    assign _1728 = ~ _1727;
    assign _130 = _91[515:515];
    always @(posedge _84) begin
        if (_82)
            _1676 <= _1675;
        else
            _1676 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1679 <= _1678;
        else
            _1679 <= _1676;
    end
    always @(posedge _84) begin
        if (_82)
            _1682 <= _1681;
        else
            _1682 <= _1679;
    end
    always @(posedge _84) begin
        if (_82)
            _1685 <= _1684;
        else
            _1685 <= _1682;
    end
    always @(posedge _84) begin
        if (_82)
            _1688 <= _1687;
        else
            _1688 <= _1685;
    end
    always @(posedge _84) begin
        if (_82)
            _1691 <= _1690;
        else
            _1691 <= _1688;
    end
    always @(posedge _84) begin
        if (_82)
            _1694 <= _1693;
        else
            _1694 <= _1691;
    end
    always @(posedge _84) begin
        if (_82)
            _1697 <= _1696;
        else
            _1697 <= _1694;
    end
    always @(posedge _84) begin
        if (_82)
            _1700 <= _1699;
        else
            _1700 <= _1697;
    end
    assign _1729 = _1700 & _1728;
    assign _102 = _91[522:522];
    always @(posedge _84) begin
        if (_82)
            _105 <= _104;
        else
            _105 <= _102;
    end
    always @(posedge _84) begin
        if (_82)
            _108 <= _107;
        else
            _108 <= _105;
    end
    always @(posedge _84) begin
        if (_82)
            _111 <= _110;
        else
            _111 <= _108;
    end
    always @(posedge _84) begin
        if (_82)
            _114 <= _113;
        else
            _114 <= _111;
    end
    always @(posedge _84) begin
        if (_82)
            _117 <= _116;
        else
            _117 <= _114;
    end
    always @(posedge _84) begin
        if (_82)
            _120 <= _119;
        else
            _120 <= _117;
    end
    always @(posedge _84) begin
        if (_82)
            _123 <= _122;
        else
            _123 <= _120;
    end
    always @(posedge _84) begin
        if (_82)
            _126 <= _125;
        else
            _126 <= _123;
    end
    always @(posedge _84) begin
        if (_82)
            _129 <= _128;
        else
            _129 <= _126;
    end
    assign _1730 = _129 & _1729;
    assign write_enable_94 = _1730 & PHASE_22;
    assign _1735 = write_enable_94 | read_enable_78;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_46
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1735), .regcea(vdd), .wea(write_enable_94), .addra(address_94), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_85), .regceb(vdd), .web(write_enable_85), .addrb(address_85), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1742[131:131]), .sbiterrb(_1742[130:130]), .doutb(_1742[129:66]), .dbiterra(_1742[65:65]), .sbiterra(_1742[64:64]), .douta(_1742[63:0]) );
    assign _1743 = _1742[63:0];
    assign _72 = flip;
    assign _1673 = ~ PHASE_22;
    assign _73 = _1673;
    always @(posedge _84) begin
        if (_82)
            PHASE_22 <= _1671;
        else
            if (_72)
                PHASE_22 <= _73;
    end
    assign _1755 = PHASE_22 ? _1754 : _1743;
    assign _76 = first_4step_pass;
    assign _78 = first_iter;
    assign _80 = start;
    assign _82 = clear;
    assign _84 = clock;
    ctrl
        ctrl
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .first_4step_pass(_76), .flip(_91[523:523]), .read_write_enable(_91[522:522]), .index(_91[521:518]), .valid(_91[517:517]), .twiddle_stage(_91[516:516]), .last_stage(_91[515:515]), .first_stage(_91[514:514]), .start_twiddles(_91[513:513]), .omegas6(_91[512:449]), .omegas5(_91[448:385]), .omegas4(_91[384:321]), .omegas3(_91[320:257]), .omegas2(_91[256:193]), .omegas1(_91[192:129]), .omegas0(_91[128:65]), .addr2(_91[64:53]), .addr1(_91[52:41]), .m(_91[40:29]), .k(_91[28:17]), .j(_91[16:5]), .i(_91[4:1]), .done_(_91[0:0]) );
    assign _1756 = _91[0:0];

    /* aliases */
    assign data_0 = data;
    assign data_2 = data_1;
    assign data_4 = data_3;
    assign data_5 = data_3;
    assign data_6 = data_3;
    assign data_8 = data_7;
    assign data_9 = data_7;
    assign data_10 = data_7;
    assign data_12 = data_11;
    assign data_14 = data_13;
    assign data_16 = data_15;
    assign data_17 = data_15;
    assign data_18 = data_15;
    assign data_20 = data_19;
    assign data_21 = data_19;
    assign data_22 = data_19;
    assign data_24 = data_23;
    assign data_26 = data_25;
    assign data_28 = data_27;
    assign data_29 = data_27;
    assign data_30 = data_27;
    assign data_32 = data_31;
    assign data_33 = data_31;
    assign data_34 = data_31;
    assign data_36 = data_35;
    assign data_38 = data_37;
    assign data_40 = data_39;
    assign data_41 = data_39;
    assign data_42 = data_39;
    assign data_44 = data_43;
    assign data_45 = data_43;
    assign data_46 = data_43;
    assign data_48 = data_47;
    assign data_50 = data_49;
    assign data_52 = data_51;
    assign data_53 = data_51;
    assign data_54 = data_51;
    assign data_56 = data_55;
    assign data_57 = data_55;
    assign data_58 = data_55;
    assign data_60 = data_59;
    assign data_62 = data_61;
    assign data_64 = data_63;
    assign data_65 = data_63;
    assign data_66 = data_63;
    assign data_68 = data_67;
    assign data_69 = data_67;
    assign data_70 = data_67;
    assign data_72 = data_71;
    assign data_74 = data_73;
    assign data_76 = data_75;
    assign data_77 = data_75;
    assign data_78 = data_75;
    assign data_80 = data_79;
    assign data_81 = data_79;
    assign data_82 = data_79;
    assign data_84 = data_83;
    assign data_86 = data_85;
    assign data_88 = data_87;
    assign data_89 = data_87;
    assign data_90 = data_87;
    assign data_92 = data_91;
    assign data_93 = data_91;
    assign data_94 = data_91;

    /* output assignments */
    assign done_ = _1756;
    assign rd_q0 = _1755;
    assign rd_q1 = _1559;
    assign rd_q2 = _1363;
    assign rd_q3 = _1167;
    assign rd_q4 = _971;
    assign rd_q5 = _775;
    assign rd_q6 = _579;
    assign rd_q7 = _383;

endmodule
module dp_23 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1011011110011011001100001001011100001010101001010000110000111110;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0011110101010110000000001101011100010100100101111100001010111100;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0101001110010000111001101101001110111101111110001100111010111111;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0110100110010111111010001101100011001001101111010100100000100101;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0000000110011111011011110111001101111001110110010011010011110001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0000101011001010001100100100101101011011001100100000011011011100;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0010101111111100010110000001100000101010110111101101100011110100;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_24 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1000001101101101010001010010111001000010111000101011100011100110;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1000101101111010111110100101101000010010011111110000010100011000;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1010011100000000010110100110101110100011001101101100100000100000;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0001011111010001110111110010100111110100110100010110100100111010;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1011001001111110010011100100101001101101101011111111101111011111;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0001100100000101011100000100110001000100110010001101110010111010;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0001011011011100101011001111000010100111110000010001101011100101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_25 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0010011101101111101110111100010110111100100101100101100000101110;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0110101010010110110001001110100010101101100101010001110111001100;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1101101101101101001101011001011000101010101101001100100010000110;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0110010010111101011010101001111010001000110111100110011111100000;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0010111110010100110000110000001100100101110011011100011011100111;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1000011011100101001000010011100100111101111001011101100010110100;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0011101010000111001111101001111000100100000111000010101101000010;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_26 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1000110100110000010001100011010110011011111001000111010101101011;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1111101101011111000100111011001000110101001100000101010001101001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1010010010110110101001100110111001101110101111010101100100111011;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0001001000111000010111110001101011011001000001111111010110000000;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1101101111000101111100101101101010110110001111000100011100110101;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0000000010100111001011000000010010100111011101011111110001111000;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0111110100110000011011110001001011110110100001101100011000110001;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_27 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1001001111001111100100101110011001000010100110100100110010010011;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1011011110011011001100001001011100001010101001010000110000111110;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1000000000010101010101101101000101010110000010111110001110111000;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0001011010011001110010100011110011001100000000011000111101010101;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0110001110111000011110101101110010111010001011110110000001100110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0100000001000101111010011110100001010111011001101011110100011101;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0000110110101000001001111111111011110100101101110111101011101101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_28 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1000000001011001111011101010000100001100000100010111011111000001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0000100110010111110010100100111100001101011111100110010000100111;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0111001011101001100010001000101100101010000111001111110010110110;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1110011011001110001111101000111100010010100010010100000110001111;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1011100001110110000110110001110011000110001011011000011111001001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0111011001011011100010101110000100110011001100001000011000011111;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1100110001010101111010011100111000000001100110010011100111110110;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_29 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0011110101010010010000101110111110001011011110110110010010111001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1010101100000000110010110011010110110001111111010100000010011110;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1000101101111010111110100101101000010010011111110000010100011000;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0101001110010000111001101101001110111101111110001100111010111111;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0100000110110111010100110011011100010101000101100000000101100101;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0101100000001101011100101110110101101100101000101100101011001111;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1101100000000001010001101110001110101111011110010110111001001011;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_30 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1011101101111110011110010101110001010010110000101001000010110101;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0011000010001100001100011100100111111111000000110100110000111001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1010111001110111011101101100110101111000100111010101001011000101;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1001000110010011001111101000110110101010110010001101001001001111;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0001100001100011000110101001001001010000010111000111101001001011;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1101101111001011010111001011111000101000101010100101110101010110;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1011100001101011010010000000101111101110010111111001010100001101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module parallel_cores_2 (
    wr_d7,
    wr_d6,
    wr_d5,
    wr_d4,
    wr_d3,
    wr_d2,
    wr_d1,
    wr_d0,
    wr_addr,
    wr_en,
    rd_addr,
    rd_en,
    flip,
    first_4step_pass,
    first_iter,
    start,
    clear,
    clock,
    done_,
    rd_q0,
    rd_q1,
    rd_q2,
    rd_q3,
    rd_q4,
    rd_q5,
    rd_q6,
    rd_q7
);

    input [63:0] wr_d7;
    input [63:0] wr_d6;
    input [63:0] wr_d5;
    input [63:0] wr_d4;
    input [63:0] wr_d3;
    input [63:0] wr_d2;
    input [63:0] wr_d1;
    input [63:0] wr_d0;
    input [11:0] wr_addr;
    input [7:0] wr_en;
    input [11:0] rd_addr;
    input [7:0] rd_en;
    input flip;
    input first_4step_pass;
    input first_iter;
    input start;
    input clear;
    input clock;
    output done_;
    output [63:0] rd_q0;
    output [63:0] rd_q1;
    output [63:0] rd_q2;
    output [63:0] rd_q3;
    output [63:0] rd_q4;
    output [63:0] rd_q5;
    output [63:0] rd_q6;
    output [63:0] rd_q7;

    /* signal declarations */
    wire [11:0] address;
    wire write_enable;
    wire [11:0] address_0;
    wire _374;
    wire read_enable;
    wire _372;
    wire write_enable_0;
    wire _376;
    wire [131:0] _381;
    wire [63:0] _382;
    wire [11:0] _367 = 12'b000000000000;
    wire [11:0] address_1;
    wire _365;
    wire write_enable_1;
    wire [63:0] _279;
    wire [63:0] _278;
    wire [63:0] _280;
    wire [63:0] _276;
    wire [63:0] _275;
    wire [63:0] q1;
    wire [63:0] _281;
    wire [11:0] address_2;
    wire write_enable_2 = 1'b0;
    wire _266;
    wire read_enable_0;
    wire [11:0] address_3;
    wire _262;
    wire read_enable_1;
    wire _260;
    wire write_enable_3;
    wire _264;
    wire [131:0] _271;
    wire [63:0] _272;
    wire [63:0] data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_0;
    wire [11:0] _254 = 12'b000000000000;
    wire _252;
    wire _251;
    wire _250;
    wire _249;
    wire _248;
    wire _247;
    wire _246;
    wire _245;
    wire _244;
    wire _243;
    wire _242;
    wire _241;
    wire [11:0] _253;
    wire [11:0] address_4;
    wire write_enable_4 = 1'b0;
    wire _238;
    wire read_enable_2;
    wire [63:0] data_1;
    wire [63:0] data_2;
    wire _235;
    wire _234;
    wire _233;
    wire _232;
    wire _231;
    wire _230;
    wire _229;
    wire _228;
    wire _227;
    wire _226;
    wire _225;
    wire _224;
    wire [11:0] _236;
    wire [11:0] address_5;
    wire _221;
    wire read_enable_3;
    wire _219;
    wire write_enable_5;
    wire _223;
    wire [131:0] _258;
    wire [63:0] _259;
    wire _87 = 1'b0;
    wire _86 = 1'b0;
    wire _89;
    wire _3;
    reg PHASE;
    wire [63:0] _273;
    wire [11:0] address_6;
    wire _211;
    wire read_enable_4;
    wire write_enable_6;
    wire _213;
    wire [11:0] address_7;
    wire _206;
    wire read_enable_5;
    wire _204;
    wire write_enable_7;
    wire _208;
    wire [131:0] _216;
    wire [63:0] _217;
    wire [63:0] _295;
    wire [63:0] data_3;
    wire [63:0] data_4;
    wire [63:0] data_5;
    wire [63:0] data_6;
    wire [11:0] address_8;
    wire _169;
    wire read_enable_6;
    wire _166;
    wire _167;
    wire write_enable_8;
    wire _171;
    wire [11:0] address_9;
    wire _134;
    wire read_enable_7;
    wire _131;
    wire _132;
    wire write_enable_9;
    wire _136;
    wire [131:0] _202;
    wire [63:0] _203;
    wire _98 = 1'b0;
    wire _97 = 1'b0;
    wire _296;
    wire _5;
    reg PHASE_0;
    wire [63:0] q0;
    wire _94 = 1'b0;
    wire _93 = 1'b0;
    reg _96;
    wire [63:0] _274;
    wire [191:0] _294;
    wire [63:0] _297;
    wire [63:0] data_7;
    wire [63:0] data_8;
    wire [63:0] data_9;
    wire [63:0] data_10;
    wire [11:0] address_10;
    wire _361;
    wire _360;
    wire read_enable_8;
    wire _354 = 1'b0;
    wire _353 = 1'b0;
    wire _351 = 1'b0;
    wire _350 = 1'b0;
    wire _348 = 1'b0;
    wire _347 = 1'b0;
    wire _345 = 1'b0;
    wire _344 = 1'b0;
    wire _342 = 1'b0;
    wire _341 = 1'b0;
    wire _339 = 1'b0;
    wire _338 = 1'b0;
    wire _336 = 1'b0;
    wire _335 = 1'b0;
    wire _333 = 1'b0;
    wire _332 = 1'b0;
    wire _330 = 1'b0;
    wire _329 = 1'b0;
    reg _331;
    reg _334;
    reg _337;
    reg _340;
    reg _343;
    reg _346;
    reg _349;
    reg _352;
    reg _355;
    wire _356;
    wire _327 = 1'b0;
    wire _326 = 1'b0;
    wire _324 = 1'b0;
    wire _323 = 1'b0;
    wire _321 = 1'b0;
    wire _320 = 1'b0;
    wire _318 = 1'b0;
    wire _317 = 1'b0;
    wire _315 = 1'b0;
    wire _314 = 1'b0;
    wire _312 = 1'b0;
    wire _311 = 1'b0;
    wire _309 = 1'b0;
    wire _308 = 1'b0;
    wire _306 = 1'b0;
    wire _305 = 1'b0;
    wire _303 = 1'b0;
    wire _302 = 1'b0;
    reg _304;
    reg _307;
    reg _310;
    reg _313;
    reg _316;
    reg _319;
    reg _322;
    reg _325;
    reg _328;
    wire _357;
    wire _358;
    wire write_enable_10;
    wire _363;
    wire [131:0] _370;
    wire [63:0] _371;
    wire _299 = 1'b0;
    wire _298 = 1'b0;
    wire _301;
    wire _7;
    reg PHASE_1;
    wire [63:0] _383;
    wire [11:0] address_11;
    wire write_enable_11;
    wire [11:0] address_12;
    wire _570;
    wire read_enable_9;
    wire _568;
    wire write_enable_12;
    wire _572;
    wire [131:0] _577;
    wire [63:0] _578;
    wire [11:0] _563 = 12'b000000000000;
    wire [11:0] address_13;
    wire _561;
    wire write_enable_13;
    wire [63:0] _486;
    wire [63:0] _485;
    wire [63:0] _487;
    wire [63:0] _483;
    wire [63:0] _482;
    wire [63:0] q1_0;
    wire [63:0] _488;
    wire [11:0] address_14;
    wire write_enable_14 = 1'b0;
    wire _473;
    wire read_enable_10;
    wire [11:0] address_15;
    wire _469;
    wire read_enable_11;
    wire _467;
    wire write_enable_15;
    wire _471;
    wire [131:0] _478;
    wire [63:0] _479;
    wire [63:0] data_11 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_12;
    wire [11:0] _461 = 12'b000000000000;
    wire _459;
    wire _458;
    wire _457;
    wire _456;
    wire _455;
    wire _454;
    wire _453;
    wire _452;
    wire _451;
    wire _450;
    wire _449;
    wire _448;
    wire [11:0] _460;
    wire [11:0] address_16;
    wire write_enable_16 = 1'b0;
    wire _445;
    wire read_enable_12;
    wire [63:0] data_13;
    wire [63:0] data_14;
    wire _442;
    wire _441;
    wire _440;
    wire _439;
    wire _438;
    wire _437;
    wire _436;
    wire _435;
    wire _434;
    wire _433;
    wire _432;
    wire _431;
    wire [11:0] _443;
    wire [11:0] address_17;
    wire _428;
    wire read_enable_13;
    wire _426;
    wire write_enable_17;
    wire _430;
    wire [131:0] _465;
    wire [63:0] _466;
    wire _385 = 1'b0;
    wire _384 = 1'b0;
    wire _387;
    wire _11;
    reg PHASE_2;
    wire [63:0] _480;
    wire [11:0] address_18;
    wire _418;
    wire read_enable_14;
    wire write_enable_18;
    wire _420;
    wire [11:0] address_19;
    wire _413;
    wire read_enable_15;
    wire _411;
    wire write_enable_19;
    wire _415;
    wire [131:0] _423;
    wire [63:0] _424;
    wire [63:0] _491;
    wire [63:0] data_15;
    wire [63:0] data_16;
    wire [63:0] data_17;
    wire [63:0] data_18;
    wire [11:0] address_20;
    wire _404;
    wire read_enable_16;
    wire _401;
    wire _402;
    wire write_enable_20;
    wire _406;
    wire [11:0] address_21;
    wire _397;
    wire read_enable_17;
    wire _394;
    wire _395;
    wire write_enable_21;
    wire _399;
    wire [131:0] _409;
    wire [63:0] _410;
    wire _392 = 1'b0;
    wire _391 = 1'b0;
    wire _492;
    wire _13;
    reg PHASE_3;
    wire [63:0] q0_0;
    wire _389 = 1'b0;
    wire _388 = 1'b0;
    reg _390;
    wire [63:0] _481;
    wire [191:0] _490;
    wire [63:0] _493;
    wire [63:0] data_19;
    wire [63:0] data_20;
    wire [63:0] data_21;
    wire [63:0] data_22;
    wire [11:0] address_22;
    wire _557;
    wire _556;
    wire read_enable_18;
    wire _550 = 1'b0;
    wire _549 = 1'b0;
    wire _547 = 1'b0;
    wire _546 = 1'b0;
    wire _544 = 1'b0;
    wire _543 = 1'b0;
    wire _541 = 1'b0;
    wire _540 = 1'b0;
    wire _538 = 1'b0;
    wire _537 = 1'b0;
    wire _535 = 1'b0;
    wire _534 = 1'b0;
    wire _532 = 1'b0;
    wire _531 = 1'b0;
    wire _529 = 1'b0;
    wire _528 = 1'b0;
    wire _526 = 1'b0;
    wire _525 = 1'b0;
    reg _527;
    reg _530;
    reg _533;
    reg _536;
    reg _539;
    reg _542;
    reg _545;
    reg _548;
    reg _551;
    wire _552;
    wire _523 = 1'b0;
    wire _522 = 1'b0;
    wire _520 = 1'b0;
    wire _519 = 1'b0;
    wire _517 = 1'b0;
    wire _516 = 1'b0;
    wire _514 = 1'b0;
    wire _513 = 1'b0;
    wire _511 = 1'b0;
    wire _510 = 1'b0;
    wire _508 = 1'b0;
    wire _507 = 1'b0;
    wire _505 = 1'b0;
    wire _504 = 1'b0;
    wire _502 = 1'b0;
    wire _501 = 1'b0;
    wire _499 = 1'b0;
    wire _498 = 1'b0;
    reg _500;
    reg _503;
    reg _506;
    reg _509;
    reg _512;
    reg _515;
    reg _518;
    reg _521;
    reg _524;
    wire _553;
    wire _554;
    wire write_enable_22;
    wire _559;
    wire [131:0] _566;
    wire [63:0] _567;
    wire _495 = 1'b0;
    wire _494 = 1'b0;
    wire _497;
    wire _15;
    reg PHASE_4;
    wire [63:0] _579;
    wire [11:0] address_23;
    wire write_enable_23;
    wire [11:0] address_24;
    wire _766;
    wire read_enable_19;
    wire _764;
    wire write_enable_24;
    wire _768;
    wire [131:0] _773;
    wire [63:0] _774;
    wire [11:0] _759 = 12'b000000000000;
    wire [11:0] address_25;
    wire _757;
    wire write_enable_25;
    wire [63:0] _682;
    wire [63:0] _681;
    wire [63:0] _683;
    wire [63:0] _679;
    wire [63:0] _678;
    wire [63:0] q1_1;
    wire [63:0] _684;
    wire [11:0] address_26;
    wire write_enable_26 = 1'b0;
    wire _669;
    wire read_enable_20;
    wire [11:0] address_27;
    wire _665;
    wire read_enable_21;
    wire _663;
    wire write_enable_27;
    wire _667;
    wire [131:0] _674;
    wire [63:0] _675;
    wire [63:0] data_23 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_24;
    wire [11:0] _657 = 12'b000000000000;
    wire _655;
    wire _654;
    wire _653;
    wire _652;
    wire _651;
    wire _650;
    wire _649;
    wire _648;
    wire _647;
    wire _646;
    wire _645;
    wire _644;
    wire [11:0] _656;
    wire [11:0] address_28;
    wire write_enable_28 = 1'b0;
    wire _641;
    wire read_enable_22;
    wire [63:0] data_25;
    wire [63:0] data_26;
    wire _638;
    wire _637;
    wire _636;
    wire _635;
    wire _634;
    wire _633;
    wire _632;
    wire _631;
    wire _630;
    wire _629;
    wire _628;
    wire _627;
    wire [11:0] _639;
    wire [11:0] address_29;
    wire _624;
    wire read_enable_23;
    wire _622;
    wire write_enable_29;
    wire _626;
    wire [131:0] _661;
    wire [63:0] _662;
    wire _581 = 1'b0;
    wire _580 = 1'b0;
    wire _583;
    wire _19;
    reg PHASE_5;
    wire [63:0] _676;
    wire [11:0] address_30;
    wire _614;
    wire read_enable_24;
    wire write_enable_30;
    wire _616;
    wire [11:0] address_31;
    wire _609;
    wire read_enable_25;
    wire _607;
    wire write_enable_31;
    wire _611;
    wire [131:0] _619;
    wire [63:0] _620;
    wire [63:0] _687;
    wire [63:0] data_27;
    wire [63:0] data_28;
    wire [63:0] data_29;
    wire [63:0] data_30;
    wire [11:0] address_32;
    wire _600;
    wire read_enable_26;
    wire _597;
    wire _598;
    wire write_enable_32;
    wire _602;
    wire [11:0] address_33;
    wire _593;
    wire read_enable_27;
    wire _590;
    wire _591;
    wire write_enable_33;
    wire _595;
    wire [131:0] _605;
    wire [63:0] _606;
    wire _588 = 1'b0;
    wire _587 = 1'b0;
    wire _688;
    wire _21;
    reg PHASE_6;
    wire [63:0] q0_1;
    wire _585 = 1'b0;
    wire _584 = 1'b0;
    reg _586;
    wire [63:0] _677;
    wire [191:0] _686;
    wire [63:0] _689;
    wire [63:0] data_31;
    wire [63:0] data_32;
    wire [63:0] data_33;
    wire [63:0] data_34;
    wire [11:0] address_34;
    wire _753;
    wire _752;
    wire read_enable_28;
    wire _746 = 1'b0;
    wire _745 = 1'b0;
    wire _743 = 1'b0;
    wire _742 = 1'b0;
    wire _740 = 1'b0;
    wire _739 = 1'b0;
    wire _737 = 1'b0;
    wire _736 = 1'b0;
    wire _734 = 1'b0;
    wire _733 = 1'b0;
    wire _731 = 1'b0;
    wire _730 = 1'b0;
    wire _728 = 1'b0;
    wire _727 = 1'b0;
    wire _725 = 1'b0;
    wire _724 = 1'b0;
    wire _722 = 1'b0;
    wire _721 = 1'b0;
    reg _723;
    reg _726;
    reg _729;
    reg _732;
    reg _735;
    reg _738;
    reg _741;
    reg _744;
    reg _747;
    wire _748;
    wire _719 = 1'b0;
    wire _718 = 1'b0;
    wire _716 = 1'b0;
    wire _715 = 1'b0;
    wire _713 = 1'b0;
    wire _712 = 1'b0;
    wire _710 = 1'b0;
    wire _709 = 1'b0;
    wire _707 = 1'b0;
    wire _706 = 1'b0;
    wire _704 = 1'b0;
    wire _703 = 1'b0;
    wire _701 = 1'b0;
    wire _700 = 1'b0;
    wire _698 = 1'b0;
    wire _697 = 1'b0;
    wire _695 = 1'b0;
    wire _694 = 1'b0;
    reg _696;
    reg _699;
    reg _702;
    reg _705;
    reg _708;
    reg _711;
    reg _714;
    reg _717;
    reg _720;
    wire _749;
    wire _750;
    wire write_enable_34;
    wire _755;
    wire [131:0] _762;
    wire [63:0] _763;
    wire _691 = 1'b0;
    wire _690 = 1'b0;
    wire _693;
    wire _23;
    reg PHASE_7;
    wire [63:0] _775;
    wire [11:0] address_35;
    wire write_enable_35;
    wire [11:0] address_36;
    wire _962;
    wire read_enable_29;
    wire _960;
    wire write_enable_36;
    wire _964;
    wire [131:0] _969;
    wire [63:0] _970;
    wire [11:0] _955 = 12'b000000000000;
    wire [11:0] address_37;
    wire _953;
    wire write_enable_37;
    wire [63:0] _878;
    wire [63:0] _877;
    wire [63:0] _879;
    wire [63:0] _875;
    wire [63:0] _874;
    wire [63:0] q1_2;
    wire [63:0] _880;
    wire [11:0] address_38;
    wire write_enable_38 = 1'b0;
    wire _865;
    wire read_enable_30;
    wire [11:0] address_39;
    wire _861;
    wire read_enable_31;
    wire _859;
    wire write_enable_39;
    wire _863;
    wire [131:0] _870;
    wire [63:0] _871;
    wire [63:0] data_35 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_36;
    wire [11:0] _853 = 12'b000000000000;
    wire _851;
    wire _850;
    wire _849;
    wire _848;
    wire _847;
    wire _846;
    wire _845;
    wire _844;
    wire _843;
    wire _842;
    wire _841;
    wire _840;
    wire [11:0] _852;
    wire [11:0] address_40;
    wire write_enable_40 = 1'b0;
    wire _837;
    wire read_enable_32;
    wire [63:0] data_37;
    wire [63:0] data_38;
    wire _834;
    wire _833;
    wire _832;
    wire _831;
    wire _830;
    wire _829;
    wire _828;
    wire _827;
    wire _826;
    wire _825;
    wire _824;
    wire _823;
    wire [11:0] _835;
    wire [11:0] address_41;
    wire _820;
    wire read_enable_33;
    wire _818;
    wire write_enable_41;
    wire _822;
    wire [131:0] _857;
    wire [63:0] _858;
    wire _777 = 1'b0;
    wire _776 = 1'b0;
    wire _779;
    wire _27;
    reg PHASE_8;
    wire [63:0] _872;
    wire [11:0] address_42;
    wire _810;
    wire read_enable_34;
    wire write_enable_42;
    wire _812;
    wire [11:0] address_43;
    wire _805;
    wire read_enable_35;
    wire _803;
    wire write_enable_43;
    wire _807;
    wire [131:0] _815;
    wire [63:0] _816;
    wire [63:0] _883;
    wire [63:0] data_39;
    wire [63:0] data_40;
    wire [63:0] data_41;
    wire [63:0] data_42;
    wire [11:0] address_44;
    wire _796;
    wire read_enable_36;
    wire _793;
    wire _794;
    wire write_enable_44;
    wire _798;
    wire [11:0] address_45;
    wire _789;
    wire read_enable_37;
    wire _786;
    wire _787;
    wire write_enable_45;
    wire _791;
    wire [131:0] _801;
    wire [63:0] _802;
    wire _784 = 1'b0;
    wire _783 = 1'b0;
    wire _884;
    wire _29;
    reg PHASE_9;
    wire [63:0] q0_2;
    wire _781 = 1'b0;
    wire _780 = 1'b0;
    reg _782;
    wire [63:0] _873;
    wire [191:0] _882;
    wire [63:0] _885;
    wire [63:0] data_43;
    wire [63:0] data_44;
    wire [63:0] data_45;
    wire [63:0] data_46;
    wire [11:0] address_46;
    wire _949;
    wire _948;
    wire read_enable_38;
    wire _942 = 1'b0;
    wire _941 = 1'b0;
    wire _939 = 1'b0;
    wire _938 = 1'b0;
    wire _936 = 1'b0;
    wire _935 = 1'b0;
    wire _933 = 1'b0;
    wire _932 = 1'b0;
    wire _930 = 1'b0;
    wire _929 = 1'b0;
    wire _927 = 1'b0;
    wire _926 = 1'b0;
    wire _924 = 1'b0;
    wire _923 = 1'b0;
    wire _921 = 1'b0;
    wire _920 = 1'b0;
    wire _918 = 1'b0;
    wire _917 = 1'b0;
    reg _919;
    reg _922;
    reg _925;
    reg _928;
    reg _931;
    reg _934;
    reg _937;
    reg _940;
    reg _943;
    wire _944;
    wire _915 = 1'b0;
    wire _914 = 1'b0;
    wire _912 = 1'b0;
    wire _911 = 1'b0;
    wire _909 = 1'b0;
    wire _908 = 1'b0;
    wire _906 = 1'b0;
    wire _905 = 1'b0;
    wire _903 = 1'b0;
    wire _902 = 1'b0;
    wire _900 = 1'b0;
    wire _899 = 1'b0;
    wire _897 = 1'b0;
    wire _896 = 1'b0;
    wire _894 = 1'b0;
    wire _893 = 1'b0;
    wire _891 = 1'b0;
    wire _890 = 1'b0;
    reg _892;
    reg _895;
    reg _898;
    reg _901;
    reg _904;
    reg _907;
    reg _910;
    reg _913;
    reg _916;
    wire _945;
    wire _946;
    wire write_enable_46;
    wire _951;
    wire [131:0] _958;
    wire [63:0] _959;
    wire _887 = 1'b0;
    wire _886 = 1'b0;
    wire _889;
    wire _31;
    reg PHASE_10;
    wire [63:0] _971;
    wire [11:0] address_47;
    wire write_enable_47;
    wire [11:0] address_48;
    wire _1158;
    wire read_enable_39;
    wire _1156;
    wire write_enable_48;
    wire _1160;
    wire [131:0] _1165;
    wire [63:0] _1166;
    wire [11:0] _1151 = 12'b000000000000;
    wire [11:0] address_49;
    wire _1149;
    wire write_enable_49;
    wire [63:0] _1074;
    wire [63:0] _1073;
    wire [63:0] _1075;
    wire [63:0] _1071;
    wire [63:0] _1070;
    wire [63:0] q1_3;
    wire [63:0] _1076;
    wire [11:0] address_50;
    wire write_enable_50 = 1'b0;
    wire _1061;
    wire read_enable_40;
    wire [11:0] address_51;
    wire _1057;
    wire read_enable_41;
    wire _1055;
    wire write_enable_51;
    wire _1059;
    wire [131:0] _1066;
    wire [63:0] _1067;
    wire [63:0] data_47 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_48;
    wire [11:0] _1049 = 12'b000000000000;
    wire _1047;
    wire _1046;
    wire _1045;
    wire _1044;
    wire _1043;
    wire _1042;
    wire _1041;
    wire _1040;
    wire _1039;
    wire _1038;
    wire _1037;
    wire _1036;
    wire [11:0] _1048;
    wire [11:0] address_52;
    wire write_enable_52 = 1'b0;
    wire _1033;
    wire read_enable_42;
    wire [63:0] data_49;
    wire [63:0] data_50;
    wire _1030;
    wire _1029;
    wire _1028;
    wire _1027;
    wire _1026;
    wire _1025;
    wire _1024;
    wire _1023;
    wire _1022;
    wire _1021;
    wire _1020;
    wire _1019;
    wire [11:0] _1031;
    wire [11:0] address_53;
    wire _1016;
    wire read_enable_43;
    wire _1014;
    wire write_enable_53;
    wire _1018;
    wire [131:0] _1053;
    wire [63:0] _1054;
    wire _973 = 1'b0;
    wire _972 = 1'b0;
    wire _975;
    wire _35;
    reg PHASE_11;
    wire [63:0] _1068;
    wire [11:0] address_54;
    wire _1006;
    wire read_enable_44;
    wire write_enable_54;
    wire _1008;
    wire [11:0] address_55;
    wire _1001;
    wire read_enable_45;
    wire _999;
    wire write_enable_55;
    wire _1003;
    wire [131:0] _1011;
    wire [63:0] _1012;
    wire [63:0] _1079;
    wire [63:0] data_51;
    wire [63:0] data_52;
    wire [63:0] data_53;
    wire [63:0] data_54;
    wire [11:0] address_56;
    wire _992;
    wire read_enable_46;
    wire _989;
    wire _990;
    wire write_enable_56;
    wire _994;
    wire [11:0] address_57;
    wire _985;
    wire read_enable_47;
    wire _982;
    wire _983;
    wire write_enable_57;
    wire _987;
    wire [131:0] _997;
    wire [63:0] _998;
    wire _980 = 1'b0;
    wire _979 = 1'b0;
    wire _1080;
    wire _37;
    reg PHASE_12;
    wire [63:0] q0_3;
    wire _977 = 1'b0;
    wire _976 = 1'b0;
    reg _978;
    wire [63:0] _1069;
    wire [191:0] _1078;
    wire [63:0] _1081;
    wire [63:0] data_55;
    wire [63:0] data_56;
    wire [63:0] data_57;
    wire [63:0] data_58;
    wire [11:0] address_58;
    wire _1145;
    wire _1144;
    wire read_enable_48;
    wire _1138 = 1'b0;
    wire _1137 = 1'b0;
    wire _1135 = 1'b0;
    wire _1134 = 1'b0;
    wire _1132 = 1'b0;
    wire _1131 = 1'b0;
    wire _1129 = 1'b0;
    wire _1128 = 1'b0;
    wire _1126 = 1'b0;
    wire _1125 = 1'b0;
    wire _1123 = 1'b0;
    wire _1122 = 1'b0;
    wire _1120 = 1'b0;
    wire _1119 = 1'b0;
    wire _1117 = 1'b0;
    wire _1116 = 1'b0;
    wire _1114 = 1'b0;
    wire _1113 = 1'b0;
    reg _1115;
    reg _1118;
    reg _1121;
    reg _1124;
    reg _1127;
    reg _1130;
    reg _1133;
    reg _1136;
    reg _1139;
    wire _1140;
    wire _1111 = 1'b0;
    wire _1110 = 1'b0;
    wire _1108 = 1'b0;
    wire _1107 = 1'b0;
    wire _1105 = 1'b0;
    wire _1104 = 1'b0;
    wire _1102 = 1'b0;
    wire _1101 = 1'b0;
    wire _1099 = 1'b0;
    wire _1098 = 1'b0;
    wire _1096 = 1'b0;
    wire _1095 = 1'b0;
    wire _1093 = 1'b0;
    wire _1092 = 1'b0;
    wire _1090 = 1'b0;
    wire _1089 = 1'b0;
    wire _1087 = 1'b0;
    wire _1086 = 1'b0;
    reg _1088;
    reg _1091;
    reg _1094;
    reg _1097;
    reg _1100;
    reg _1103;
    reg _1106;
    reg _1109;
    reg _1112;
    wire _1141;
    wire _1142;
    wire write_enable_58;
    wire _1147;
    wire [131:0] _1154;
    wire [63:0] _1155;
    wire _1083 = 1'b0;
    wire _1082 = 1'b0;
    wire _1085;
    wire _39;
    reg PHASE_13;
    wire [63:0] _1167;
    wire [11:0] address_59;
    wire write_enable_59;
    wire [11:0] address_60;
    wire _1354;
    wire read_enable_49;
    wire _1352;
    wire write_enable_60;
    wire _1356;
    wire [131:0] _1361;
    wire [63:0] _1362;
    wire [11:0] _1347 = 12'b000000000000;
    wire [11:0] address_61;
    wire _1345;
    wire write_enable_61;
    wire [63:0] _1270;
    wire [63:0] _1269;
    wire [63:0] _1271;
    wire [63:0] _1267;
    wire [63:0] _1266;
    wire [63:0] q1_4;
    wire [63:0] _1272;
    wire [11:0] address_62;
    wire write_enable_62 = 1'b0;
    wire _1257;
    wire read_enable_50;
    wire [11:0] address_63;
    wire _1253;
    wire read_enable_51;
    wire _1251;
    wire write_enable_63;
    wire _1255;
    wire [131:0] _1262;
    wire [63:0] _1263;
    wire [63:0] data_59 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_60;
    wire [11:0] _1245 = 12'b000000000000;
    wire _1243;
    wire _1242;
    wire _1241;
    wire _1240;
    wire _1239;
    wire _1238;
    wire _1237;
    wire _1236;
    wire _1235;
    wire _1234;
    wire _1233;
    wire _1232;
    wire [11:0] _1244;
    wire [11:0] address_64;
    wire write_enable_64 = 1'b0;
    wire _1229;
    wire read_enable_52;
    wire [63:0] data_61;
    wire [63:0] data_62;
    wire _1226;
    wire _1225;
    wire _1224;
    wire _1223;
    wire _1222;
    wire _1221;
    wire _1220;
    wire _1219;
    wire _1218;
    wire _1217;
    wire _1216;
    wire _1215;
    wire [11:0] _1227;
    wire [11:0] address_65;
    wire _1212;
    wire read_enable_53;
    wire _1210;
    wire write_enable_65;
    wire _1214;
    wire [131:0] _1249;
    wire [63:0] _1250;
    wire _1169 = 1'b0;
    wire _1168 = 1'b0;
    wire _1171;
    wire _43;
    reg PHASE_14;
    wire [63:0] _1264;
    wire [11:0] address_66;
    wire _1202;
    wire read_enable_54;
    wire write_enable_66;
    wire _1204;
    wire [11:0] address_67;
    wire _1197;
    wire read_enable_55;
    wire _1195;
    wire write_enable_67;
    wire _1199;
    wire [131:0] _1207;
    wire [63:0] _1208;
    wire [63:0] _1275;
    wire [63:0] data_63;
    wire [63:0] data_64;
    wire [63:0] data_65;
    wire [63:0] data_66;
    wire [11:0] address_68;
    wire _1188;
    wire read_enable_56;
    wire _1185;
    wire _1186;
    wire write_enable_68;
    wire _1190;
    wire [11:0] address_69;
    wire _1181;
    wire read_enable_57;
    wire _1178;
    wire _1179;
    wire write_enable_69;
    wire _1183;
    wire [131:0] _1193;
    wire [63:0] _1194;
    wire _1176 = 1'b0;
    wire _1175 = 1'b0;
    wire _1276;
    wire _45;
    reg PHASE_15;
    wire [63:0] q0_4;
    wire _1173 = 1'b0;
    wire _1172 = 1'b0;
    reg _1174;
    wire [63:0] _1265;
    wire [191:0] _1274;
    wire [63:0] _1277;
    wire [63:0] data_67;
    wire [63:0] data_68;
    wire [63:0] data_69;
    wire [63:0] data_70;
    wire [11:0] address_70;
    wire _1341;
    wire _1340;
    wire read_enable_58;
    wire _1334 = 1'b0;
    wire _1333 = 1'b0;
    wire _1331 = 1'b0;
    wire _1330 = 1'b0;
    wire _1328 = 1'b0;
    wire _1327 = 1'b0;
    wire _1325 = 1'b0;
    wire _1324 = 1'b0;
    wire _1322 = 1'b0;
    wire _1321 = 1'b0;
    wire _1319 = 1'b0;
    wire _1318 = 1'b0;
    wire _1316 = 1'b0;
    wire _1315 = 1'b0;
    wire _1313 = 1'b0;
    wire _1312 = 1'b0;
    wire _1310 = 1'b0;
    wire _1309 = 1'b0;
    reg _1311;
    reg _1314;
    reg _1317;
    reg _1320;
    reg _1323;
    reg _1326;
    reg _1329;
    reg _1332;
    reg _1335;
    wire _1336;
    wire _1307 = 1'b0;
    wire _1306 = 1'b0;
    wire _1304 = 1'b0;
    wire _1303 = 1'b0;
    wire _1301 = 1'b0;
    wire _1300 = 1'b0;
    wire _1298 = 1'b0;
    wire _1297 = 1'b0;
    wire _1295 = 1'b0;
    wire _1294 = 1'b0;
    wire _1292 = 1'b0;
    wire _1291 = 1'b0;
    wire _1289 = 1'b0;
    wire _1288 = 1'b0;
    wire _1286 = 1'b0;
    wire _1285 = 1'b0;
    wire _1283 = 1'b0;
    wire _1282 = 1'b0;
    reg _1284;
    reg _1287;
    reg _1290;
    reg _1293;
    reg _1296;
    reg _1299;
    reg _1302;
    reg _1305;
    reg _1308;
    wire _1337;
    wire _1338;
    wire write_enable_70;
    wire _1343;
    wire [131:0] _1350;
    wire [63:0] _1351;
    wire _1279 = 1'b0;
    wire _1278 = 1'b0;
    wire _1281;
    wire _47;
    reg PHASE_16;
    wire [63:0] _1363;
    wire [11:0] address_71;
    wire write_enable_71;
    wire [11:0] address_72;
    wire _1550;
    wire read_enable_59;
    wire _1548;
    wire write_enable_72;
    wire _1552;
    wire [131:0] _1557;
    wire [63:0] _1558;
    wire [11:0] _1543 = 12'b000000000000;
    wire [11:0] address_73;
    wire _1541;
    wire write_enable_73;
    wire [63:0] _1466;
    wire [63:0] _1465;
    wire [63:0] _1467;
    wire [63:0] _1463;
    wire [63:0] _1462;
    wire [63:0] q1_5;
    wire [63:0] _1468;
    wire [11:0] address_74;
    wire write_enable_74 = 1'b0;
    wire _1453;
    wire read_enable_60;
    wire [11:0] address_75;
    wire _1449;
    wire read_enable_61;
    wire _1447;
    wire write_enable_75;
    wire _1451;
    wire [131:0] _1458;
    wire [63:0] _1459;
    wire [63:0] data_71 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_72;
    wire [11:0] _1441 = 12'b000000000000;
    wire _1439;
    wire _1438;
    wire _1437;
    wire _1436;
    wire _1435;
    wire _1434;
    wire _1433;
    wire _1432;
    wire _1431;
    wire _1430;
    wire _1429;
    wire _1428;
    wire [11:0] _1440;
    wire [11:0] address_76;
    wire write_enable_76 = 1'b0;
    wire _1425;
    wire read_enable_62;
    wire [63:0] data_73;
    wire [63:0] data_74;
    wire _1422;
    wire _1421;
    wire _1420;
    wire _1419;
    wire _1418;
    wire _1417;
    wire _1416;
    wire _1415;
    wire _1414;
    wire _1413;
    wire _1412;
    wire _1411;
    wire [11:0] _1423;
    wire [11:0] address_77;
    wire _1408;
    wire read_enable_63;
    wire _1406;
    wire write_enable_77;
    wire _1410;
    wire [131:0] _1445;
    wire [63:0] _1446;
    wire _1365 = 1'b0;
    wire _1364 = 1'b0;
    wire _1367;
    wire _51;
    reg PHASE_17;
    wire [63:0] _1460;
    wire [11:0] address_78;
    wire _1398;
    wire read_enable_64;
    wire write_enable_78;
    wire _1400;
    wire [11:0] address_79;
    wire _1393;
    wire read_enable_65;
    wire _1391;
    wire write_enable_79;
    wire _1395;
    wire [131:0] _1403;
    wire [63:0] _1404;
    wire [63:0] _1471;
    wire [63:0] data_75;
    wire [63:0] data_76;
    wire [63:0] data_77;
    wire [63:0] data_78;
    wire [11:0] address_80;
    wire _1384;
    wire read_enable_66;
    wire _1381;
    wire _1382;
    wire write_enable_80;
    wire _1386;
    wire [11:0] address_81;
    wire _1377;
    wire read_enable_67;
    wire _1374;
    wire _1375;
    wire write_enable_81;
    wire _1379;
    wire [131:0] _1389;
    wire [63:0] _1390;
    wire _1372 = 1'b0;
    wire _1371 = 1'b0;
    wire _1472;
    wire _53;
    reg PHASE_18;
    wire [63:0] q0_5;
    wire _1369 = 1'b0;
    wire _1368 = 1'b0;
    reg _1370;
    wire [63:0] _1461;
    wire [191:0] _1470;
    wire [63:0] _1473;
    wire [63:0] data_79;
    wire [63:0] data_80;
    wire [63:0] data_81;
    wire [63:0] data_82;
    wire [11:0] address_82;
    wire _1537;
    wire _1536;
    wire read_enable_68;
    wire _1530 = 1'b0;
    wire _1529 = 1'b0;
    wire _1527 = 1'b0;
    wire _1526 = 1'b0;
    wire _1524 = 1'b0;
    wire _1523 = 1'b0;
    wire _1521 = 1'b0;
    wire _1520 = 1'b0;
    wire _1518 = 1'b0;
    wire _1517 = 1'b0;
    wire _1515 = 1'b0;
    wire _1514 = 1'b0;
    wire _1512 = 1'b0;
    wire _1511 = 1'b0;
    wire _1509 = 1'b0;
    wire _1508 = 1'b0;
    wire _1506 = 1'b0;
    wire _1505 = 1'b0;
    reg _1507;
    reg _1510;
    reg _1513;
    reg _1516;
    reg _1519;
    reg _1522;
    reg _1525;
    reg _1528;
    reg _1531;
    wire _1532;
    wire _1503 = 1'b0;
    wire _1502 = 1'b0;
    wire _1500 = 1'b0;
    wire _1499 = 1'b0;
    wire _1497 = 1'b0;
    wire _1496 = 1'b0;
    wire _1494 = 1'b0;
    wire _1493 = 1'b0;
    wire _1491 = 1'b0;
    wire _1490 = 1'b0;
    wire _1488 = 1'b0;
    wire _1487 = 1'b0;
    wire _1485 = 1'b0;
    wire _1484 = 1'b0;
    wire _1482 = 1'b0;
    wire _1481 = 1'b0;
    wire _1479 = 1'b0;
    wire _1478 = 1'b0;
    reg _1480;
    reg _1483;
    reg _1486;
    reg _1489;
    reg _1492;
    reg _1495;
    reg _1498;
    reg _1501;
    reg _1504;
    wire _1533;
    wire _1534;
    wire write_enable_82;
    wire _1539;
    wire [131:0] _1546;
    wire [63:0] _1547;
    wire _1475 = 1'b0;
    wire _1474 = 1'b0;
    wire _1477;
    wire _55;
    reg PHASE_19;
    wire [63:0] _1559;
    wire [11:0] address_83;
    wire write_enable_83;
    wire [11:0] address_84;
    wire _1746;
    wire read_enable_69;
    wire _1744;
    wire write_enable_84;
    wire _1748;
    wire [131:0] _1753;
    wire [63:0] _1754;
    wire [11:0] _1739 = 12'b000000000000;
    wire [11:0] address_85;
    wire _1737;
    wire write_enable_85;
    wire [3:0] _292;
    wire _291;
    wire _289;
    wire [63:0] _288;
    wire [63:0] _287;
    wire [63:0] _286;
    wire [63:0] _285;
    wire [63:0] _284;
    wire [63:0] _283;
    wire [63:0] _282;
    wire [63:0] _1662;
    wire [63:0] _1661;
    wire [63:0] _1663;
    wire [63:0] _1659;
    wire [63:0] _1658;
    wire [63:0] q1_6;
    wire [63:0] _1664;
    wire [11:0] address_86;
    wire write_enable_86 = 1'b0;
    wire _1649;
    wire read_enable_70;
    wire [11:0] address_87;
    wire _1645;
    wire read_enable_71;
    wire _1643;
    wire write_enable_87;
    wire _1647;
    wire [131:0] _1654;
    wire [63:0] _1655;
    wire [63:0] data_83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_84;
    wire [11:0] _1637 = 12'b000000000000;
    wire _1635;
    wire _1634;
    wire _1633;
    wire _1632;
    wire _1631;
    wire _1630;
    wire _1629;
    wire _1628;
    wire _1627;
    wire _1626;
    wire _1625;
    wire _1624;
    wire [11:0] _1636;
    wire [11:0] address_88;
    wire write_enable_88 = 1'b0;
    wire _1621;
    wire read_enable_72;
    wire [63:0] data_85;
    wire [63:0] data_86;
    wire [11:0] _60;
    wire _1618;
    wire _1617;
    wire _1616;
    wire _1615;
    wire _1614;
    wire _1613;
    wire _1612;
    wire _1611;
    wire _1610;
    wire _1609;
    wire _1608;
    wire _1607;
    wire [11:0] _1619;
    wire [11:0] address_89;
    wire _1604;
    wire read_enable_73;
    wire [7:0] _62;
    wire _1602;
    wire write_enable_89;
    wire _1606;
    wire [131:0] _1641;
    wire [63:0] _1642;
    wire _1561 = 1'b0;
    wire _1560 = 1'b0;
    wire _1563;
    wire _63;
    reg PHASE_20;
    wire [63:0] _1656;
    wire [11:0] address_90;
    wire _1594;
    wire read_enable_74;
    wire write_enable_90;
    wire _1596;
    wire [11:0] address_91;
    wire _1589;
    wire read_enable_75;
    wire _1587;
    wire write_enable_91;
    wire _1591;
    wire [131:0] _1599;
    wire [63:0] _1600;
    wire [63:0] _1667;
    wire [63:0] data_87;
    wire [63:0] data_88;
    wire [63:0] data_89;
    wire [63:0] data_90;
    wire [11:0] _198 = 12'b000000000000;
    wire [11:0] _197 = 12'b000000000000;
    wire [11:0] _195 = 12'b000000000000;
    wire [11:0] _194 = 12'b000000000000;
    wire [11:0] _192 = 12'b000000000000;
    wire [11:0] _191 = 12'b000000000000;
    wire [11:0] _189 = 12'b000000000000;
    wire [11:0] _188 = 12'b000000000000;
    wire [11:0] _186 = 12'b000000000000;
    wire [11:0] _185 = 12'b000000000000;
    wire [11:0] _183 = 12'b000000000000;
    wire [11:0] _182 = 12'b000000000000;
    wire [11:0] _180 = 12'b000000000000;
    wire [11:0] _179 = 12'b000000000000;
    wire [11:0] _177 = 12'b000000000000;
    wire [11:0] _176 = 12'b000000000000;
    wire [11:0] _174 = 12'b000000000000;
    wire [11:0] _173 = 12'b000000000000;
    reg [11:0] _175;
    reg [11:0] _178;
    reg [11:0] _181;
    reg [11:0] _184;
    reg [11:0] _187;
    reg [11:0] _190;
    reg [11:0] _193;
    reg [11:0] _196;
    reg [11:0] _199;
    wire [11:0] _172;
    wire [11:0] address_92;
    wire _1580;
    wire read_enable_76;
    wire _1577;
    wire _1578;
    wire write_enable_92;
    wire _1582;
    wire [11:0] address_93;
    wire _1573;
    wire read_enable_77;
    wire _1570;
    wire _1571;
    wire write_enable_93;
    wire _1575;
    wire [131:0] _1585;
    wire [63:0] _1586;
    wire _99;
    wire _1568 = 1'b0;
    wire _1567 = 1'b0;
    wire _1668;
    wire _65;
    reg PHASE_21;
    wire [63:0] q0_6;
    wire _1565 = 1'b0;
    wire _1564 = 1'b0;
    wire _92;
    reg _1566;
    wire [63:0] _1657;
    wire [191:0] _1666;
    wire [63:0] _1669;
    wire [63:0] data_91;
    wire [63:0] data_92;
    wire [63:0] data_93;
    wire [63:0] data_94;
    wire [11:0] _163 = 12'b000000000000;
    wire [11:0] _162 = 12'b000000000000;
    wire [11:0] _160 = 12'b000000000000;
    wire [11:0] _159 = 12'b000000000000;
    wire [11:0] _157 = 12'b000000000000;
    wire [11:0] _156 = 12'b000000000000;
    wire [11:0] _154 = 12'b000000000000;
    wire [11:0] _153 = 12'b000000000000;
    wire [11:0] _151 = 12'b000000000000;
    wire [11:0] _150 = 12'b000000000000;
    wire [11:0] _148 = 12'b000000000000;
    wire [11:0] _147 = 12'b000000000000;
    wire [11:0] _145 = 12'b000000000000;
    wire [11:0] _144 = 12'b000000000000;
    wire [11:0] _142 = 12'b000000000000;
    wire [11:0] _141 = 12'b000000000000;
    wire [11:0] _139 = 12'b000000000000;
    wire [11:0] _138 = 12'b000000000000;
    wire [11:0] _137;
    reg [11:0] _140;
    reg [11:0] _143;
    reg [11:0] _146;
    reg [11:0] _149;
    reg [11:0] _152;
    reg [11:0] _155;
    reg [11:0] _158;
    reg [11:0] _161;
    reg [11:0] _164;
    wire [11:0] _68;
    wire [11:0] address_94;
    wire _1733;
    wire [7:0] _70;
    wire _1732;
    wire read_enable_78;
    wire _1726 = 1'b0;
    wire _1725 = 1'b0;
    wire _1723 = 1'b0;
    wire _1722 = 1'b0;
    wire _1720 = 1'b0;
    wire _1719 = 1'b0;
    wire _1717 = 1'b0;
    wire _1716 = 1'b0;
    wire _1714 = 1'b0;
    wire _1713 = 1'b0;
    wire _1711 = 1'b0;
    wire _1710 = 1'b0;
    wire _1708 = 1'b0;
    wire _1707 = 1'b0;
    wire _1705 = 1'b0;
    wire _1704 = 1'b0;
    wire _1702 = 1'b0;
    wire _1701 = 1'b0;
    wire _290;
    reg _1703;
    reg _1706;
    reg _1709;
    reg _1712;
    reg _1715;
    reg _1718;
    reg _1721;
    reg _1724;
    reg _1727;
    wire _1728;
    wire _1699 = 1'b0;
    wire _1698 = 1'b0;
    wire _1696 = 1'b0;
    wire _1695 = 1'b0;
    wire _1693 = 1'b0;
    wire _1692 = 1'b0;
    wire _1690 = 1'b0;
    wire _1689 = 1'b0;
    wire _1687 = 1'b0;
    wire _1686 = 1'b0;
    wire _1684 = 1'b0;
    wire _1683 = 1'b0;
    wire _1681 = 1'b0;
    wire _1680 = 1'b0;
    wire _1678 = 1'b0;
    wire _1677 = 1'b0;
    wire _1675 = 1'b0;
    wire _1674 = 1'b0;
    wire _130;
    reg _1676;
    reg _1679;
    reg _1682;
    reg _1685;
    reg _1688;
    reg _1691;
    reg _1694;
    reg _1697;
    reg _1700;
    wire _1729;
    wire _128 = 1'b0;
    wire _127 = 1'b0;
    wire _125 = 1'b0;
    wire _124 = 1'b0;
    wire _122 = 1'b0;
    wire _121 = 1'b0;
    wire _119 = 1'b0;
    wire _118 = 1'b0;
    wire _116 = 1'b0;
    wire _115 = 1'b0;
    wire _113 = 1'b0;
    wire _112 = 1'b0;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire vdd = 1'b1;
    wire _104 = 1'b0;
    wire _103 = 1'b0;
    wire _102;
    reg _105;
    reg _108;
    reg _111;
    reg _114;
    reg _117;
    reg _120;
    reg _123;
    reg _126;
    reg _129;
    wire _1730;
    wire write_enable_94;
    wire _1735;
    wire gnd = 1'b0;
    wire [131:0] _1742;
    wire [63:0] _1743;
    wire _72;
    wire _1671 = 1'b0;
    wire _1670 = 1'b0;
    wire _1673;
    wire _73;
    reg PHASE_22;
    wire [63:0] _1755;
    wire _76;
    wire _78;
    wire _80;
    wire _82;
    wire _84;
    wire [523:0] _91;
    wire _1756;

    /* logic */
    assign address = _372 ? _199 : _367;
    assign write_enable = _365 & _372;
    assign address_0 = _372 ? _164 : _68;
    assign _374 = ~ _372;
    assign read_enable = _360 & _374;
    assign _372 = ~ PHASE_1;
    assign write_enable_0 = _358 & _372;
    assign _376 = write_enable_0 | read_enable;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_376), .regcea(vdd), .wea(write_enable_0), .addra(address_0), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable), .regceb(vdd), .web(write_enable), .addrb(address), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_381[131:131]), .sbiterrb(_381[130:130]), .doutb(_381[129:66]), .dbiterra(_381[65:65]), .sbiterra(_381[64:64]), .douta(_381[63:0]) );
    assign _382 = _381[63:0];
    assign address_1 = PHASE_1 ? _199 : _367;
    assign _365 = _129 & _328;
    assign write_enable_1 = _365 & PHASE_1;
    assign _279 = _271[129:66];
    assign _278 = _258[129:66];
    assign _280 = PHASE ? _279 : _278;
    assign _276 = _216[129:66];
    assign _275 = _202[129:66];
    assign q1 = PHASE_0 ? _276 : _275;
    assign _281 = _96 ? _280 : q1;
    assign address_2 = _260 ? _254 : _253;
    assign _266 = ~ _260;
    assign read_enable_0 = _102 & _266;
    assign address_3 = _260 ? _60 : _236;
    assign _262 = ~ _260;
    assign read_enable_1 = _102 & _262;
    assign _260 = ~ PHASE;
    assign write_enable_3 = _219 & _260;
    assign _264 = write_enable_3 | read_enable_1;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_0
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_264), .regcea(vdd), .wea(write_enable_3), .addra(address_3), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_0), .regceb(vdd), .web(write_enable_2), .addrb(address_2), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_271[131:131]), .sbiterrb(_271[130:130]), .doutb(_271[129:66]), .dbiterra(_271[65:65]), .sbiterra(_271[64:64]), .douta(_271[63:0]) );
    assign _272 = _271[63:0];
    assign _252 = _172[11:11];
    assign _251 = _172[10:10];
    assign _250 = _172[9:9];
    assign _249 = _172[8:8];
    assign _248 = _172[7:7];
    assign _247 = _172[6:6];
    assign _246 = _172[5:5];
    assign _245 = _172[4:4];
    assign _244 = _172[3:3];
    assign _243 = _172[2:2];
    assign _242 = _172[1:1];
    assign _241 = _172[0:0];
    assign _253 = { _241, _242, _243, _244, _245, _246, _247, _248, _249, _250, _251, _252 };
    assign address_4 = PHASE ? _254 : _253;
    assign _238 = ~ PHASE;
    assign read_enable_2 = _102 & _238;
    assign data_1 = wr_d7;
    assign _235 = _137[11:11];
    assign _234 = _137[10:10];
    assign _233 = _137[9:9];
    assign _232 = _137[8:8];
    assign _231 = _137[7:7];
    assign _230 = _137[6:6];
    assign _229 = _137[5:5];
    assign _228 = _137[4:4];
    assign _227 = _137[3:3];
    assign _226 = _137[2:2];
    assign _225 = _137[1:1];
    assign _224 = _137[0:0];
    assign _236 = { _224, _225, _226, _227, _228, _229, _230, _231, _232, _233, _234, _235 };
    assign address_5 = PHASE ? _60 : _236;
    assign _221 = ~ PHASE;
    assign read_enable_3 = _102 & _221;
    assign _219 = _62[7:7];
    assign write_enable_5 = _219 & PHASE;
    assign _223 = write_enable_5 | read_enable_3;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_1
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_223), .regcea(vdd), .wea(write_enable_5), .addra(address_5), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_2), .regceb(vdd), .web(write_enable_4), .addrb(address_4), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_258[131:131]), .sbiterrb(_258[130:130]), .doutb(_258[129:66]), .dbiterra(_258[65:65]), .sbiterra(_258[64:64]), .douta(_258[63:0]) );
    assign _259 = _258[63:0];
    assign _89 = ~ PHASE;
    assign _3 = _89;
    always @(posedge _84) begin
        if (_82)
            PHASE <= _87;
        else
            if (_72)
                PHASE <= _3;
    end
    assign _273 = PHASE ? _272 : _259;
    assign address_6 = _204 ? _199 : _172;
    assign _211 = ~ _204;
    assign read_enable_4 = _102 & _211;
    assign write_enable_6 = _167 & _204;
    assign _213 = write_enable_6 | read_enable_4;
    assign address_7 = _204 ? _164 : _137;
    assign _206 = ~ _204;
    assign read_enable_5 = _102 & _206;
    assign _204 = ~ PHASE_0;
    assign write_enable_7 = _132 & _204;
    assign _208 = write_enable_7 | read_enable_5;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_2
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_208), .regcea(vdd), .wea(write_enable_7), .addra(address_7), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_213), .regceb(vdd), .web(write_enable_6), .addrb(address_6), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_216[131:131]), .sbiterrb(_216[130:130]), .doutb(_216[129:66]), .dbiterra(_216[65:65]), .sbiterra(_216[64:64]), .douta(_216[63:0]) );
    assign _217 = _216[63:0];
    assign _295 = _294[127:64];
    assign data_3 = _295;
    assign address_8 = PHASE_0 ? _199 : _172;
    assign _169 = ~ PHASE_0;
    assign read_enable_6 = _102 & _169;
    assign _166 = ~ _130;
    assign _167 = _129 & _166;
    assign write_enable_8 = _167 & PHASE_0;
    assign _171 = write_enable_8 | read_enable_6;
    assign address_9 = PHASE_0 ? _164 : _137;
    assign _134 = ~ PHASE_0;
    assign read_enable_7 = _102 & _134;
    assign _131 = ~ _130;
    assign _132 = _129 & _131;
    assign write_enable_9 = _132 & PHASE_0;
    assign _136 = write_enable_9 | read_enable_7;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_3
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_136), .regcea(vdd), .wea(write_enable_9), .addra(address_9), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_171), .regceb(vdd), .web(write_enable_8), .addrb(address_8), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_202[131:131]), .sbiterrb(_202[130:130]), .doutb(_202[129:66]), .dbiterra(_202[65:65]), .sbiterra(_202[64:64]), .douta(_202[63:0]) );
    assign _203 = _202[63:0];
    assign _296 = ~ PHASE_0;
    assign _5 = _296;
    always @(posedge _84) begin
        if (_82)
            PHASE_0 <= _98;
        else
            if (_99)
                PHASE_0 <= _5;
    end
    assign q0 = PHASE_0 ? _217 : _203;
    always @(posedge _84) begin
        if (_82)
            _96 <= _94;
        else
            _96 <= _92;
    end
    assign _274 = _96 ? _273 : q0;
    dp_30
        dp_6
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_274), .d2(_281), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_294[191:128]), .q2(_294[127:64]), .q1(_294[63:0]) );
    assign _297 = _294[63:0];
    assign data_7 = _297;
    assign address_10 = PHASE_1 ? _164 : _68;
    assign _361 = ~ PHASE_1;
    assign _360 = _70[7:7];
    assign read_enable_8 = _360 & _361;
    always @(posedge _84) begin
        if (_82)
            _331 <= _330;
        else
            _331 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _334 <= _333;
        else
            _334 <= _331;
    end
    always @(posedge _84) begin
        if (_82)
            _337 <= _336;
        else
            _337 <= _334;
    end
    always @(posedge _84) begin
        if (_82)
            _340 <= _339;
        else
            _340 <= _337;
    end
    always @(posedge _84) begin
        if (_82)
            _343 <= _342;
        else
            _343 <= _340;
    end
    always @(posedge _84) begin
        if (_82)
            _346 <= _345;
        else
            _346 <= _343;
    end
    always @(posedge _84) begin
        if (_82)
            _349 <= _348;
        else
            _349 <= _346;
    end
    always @(posedge _84) begin
        if (_82)
            _352 <= _351;
        else
            _352 <= _349;
    end
    always @(posedge _84) begin
        if (_82)
            _355 <= _354;
        else
            _355 <= _352;
    end
    assign _356 = ~ _355;
    always @(posedge _84) begin
        if (_82)
            _304 <= _303;
        else
            _304 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _307 <= _306;
        else
            _307 <= _304;
    end
    always @(posedge _84) begin
        if (_82)
            _310 <= _309;
        else
            _310 <= _307;
    end
    always @(posedge _84) begin
        if (_82)
            _313 <= _312;
        else
            _313 <= _310;
    end
    always @(posedge _84) begin
        if (_82)
            _316 <= _315;
        else
            _316 <= _313;
    end
    always @(posedge _84) begin
        if (_82)
            _319 <= _318;
        else
            _319 <= _316;
    end
    always @(posedge _84) begin
        if (_82)
            _322 <= _321;
        else
            _322 <= _319;
    end
    always @(posedge _84) begin
        if (_82)
            _325 <= _324;
        else
            _325 <= _322;
    end
    always @(posedge _84) begin
        if (_82)
            _328 <= _327;
        else
            _328 <= _325;
    end
    assign _357 = _328 & _356;
    assign _358 = _129 & _357;
    assign write_enable_10 = _358 & PHASE_1;
    assign _363 = write_enable_10 | read_enable_8;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_4
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_363), .regcea(vdd), .wea(write_enable_10), .addra(address_10), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_1), .regceb(vdd), .web(write_enable_1), .addrb(address_1), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_370[131:131]), .sbiterrb(_370[130:130]), .doutb(_370[129:66]), .dbiterra(_370[65:65]), .sbiterra(_370[64:64]), .douta(_370[63:0]) );
    assign _371 = _370[63:0];
    assign _301 = ~ PHASE_1;
    assign _7 = _301;
    always @(posedge _84) begin
        if (_82)
            PHASE_1 <= _299;
        else
            if (_72)
                PHASE_1 <= _7;
    end
    assign _383 = PHASE_1 ? _382 : _371;
    assign address_11 = _568 ? _199 : _563;
    assign write_enable_11 = _561 & _568;
    assign address_12 = _568 ? _164 : _68;
    assign _570 = ~ _568;
    assign read_enable_9 = _556 & _570;
    assign _568 = ~ PHASE_4;
    assign write_enable_12 = _554 & _568;
    assign _572 = write_enable_12 | read_enable_9;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_5
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_572), .regcea(vdd), .wea(write_enable_12), .addra(address_12), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_11), .regceb(vdd), .web(write_enable_11), .addrb(address_11), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_577[131:131]), .sbiterrb(_577[130:130]), .doutb(_577[129:66]), .dbiterra(_577[65:65]), .sbiterra(_577[64:64]), .douta(_577[63:0]) );
    assign _578 = _577[63:0];
    assign address_13 = PHASE_4 ? _199 : _563;
    assign _561 = _129 & _524;
    assign write_enable_13 = _561 & PHASE_4;
    assign _486 = _478[129:66];
    assign _485 = _465[129:66];
    assign _487 = PHASE_2 ? _486 : _485;
    assign _483 = _423[129:66];
    assign _482 = _409[129:66];
    assign q1_0 = PHASE_3 ? _483 : _482;
    assign _488 = _390 ? _487 : q1_0;
    assign address_14 = _467 ? _461 : _460;
    assign _473 = ~ _467;
    assign read_enable_10 = _102 & _473;
    assign address_15 = _467 ? _60 : _443;
    assign _469 = ~ _467;
    assign read_enable_11 = _102 & _469;
    assign _467 = ~ PHASE_2;
    assign write_enable_15 = _426 & _467;
    assign _471 = write_enable_15 | read_enable_11;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_6
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_471), .regcea(vdd), .wea(write_enable_15), .addra(address_15), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_10), .regceb(vdd), .web(write_enable_14), .addrb(address_14), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_478[131:131]), .sbiterrb(_478[130:130]), .doutb(_478[129:66]), .dbiterra(_478[65:65]), .sbiterra(_478[64:64]), .douta(_478[63:0]) );
    assign _479 = _478[63:0];
    assign _459 = _172[11:11];
    assign _458 = _172[10:10];
    assign _457 = _172[9:9];
    assign _456 = _172[8:8];
    assign _455 = _172[7:7];
    assign _454 = _172[6:6];
    assign _453 = _172[5:5];
    assign _452 = _172[4:4];
    assign _451 = _172[3:3];
    assign _450 = _172[2:2];
    assign _449 = _172[1:1];
    assign _448 = _172[0:0];
    assign _460 = { _448, _449, _450, _451, _452, _453, _454, _455, _456, _457, _458, _459 };
    assign address_16 = PHASE_2 ? _461 : _460;
    assign _445 = ~ PHASE_2;
    assign read_enable_12 = _102 & _445;
    assign data_13 = wr_d6;
    assign _442 = _137[11:11];
    assign _441 = _137[10:10];
    assign _440 = _137[9:9];
    assign _439 = _137[8:8];
    assign _438 = _137[7:7];
    assign _437 = _137[6:6];
    assign _436 = _137[5:5];
    assign _435 = _137[4:4];
    assign _434 = _137[3:3];
    assign _433 = _137[2:2];
    assign _432 = _137[1:1];
    assign _431 = _137[0:0];
    assign _443 = { _431, _432, _433, _434, _435, _436, _437, _438, _439, _440, _441, _442 };
    assign address_17 = PHASE_2 ? _60 : _443;
    assign _428 = ~ PHASE_2;
    assign read_enable_13 = _102 & _428;
    assign _426 = _62[6:6];
    assign write_enable_17 = _426 & PHASE_2;
    assign _430 = write_enable_17 | read_enable_13;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_7
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_430), .regcea(vdd), .wea(write_enable_17), .addra(address_17), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_12), .regceb(vdd), .web(write_enable_16), .addrb(address_16), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_465[131:131]), .sbiterrb(_465[130:130]), .doutb(_465[129:66]), .dbiterra(_465[65:65]), .sbiterra(_465[64:64]), .douta(_465[63:0]) );
    assign _466 = _465[63:0];
    assign _387 = ~ PHASE_2;
    assign _11 = _387;
    always @(posedge _84) begin
        if (_82)
            PHASE_2 <= _385;
        else
            if (_72)
                PHASE_2 <= _11;
    end
    assign _480 = PHASE_2 ? _479 : _466;
    assign address_18 = _411 ? _199 : _172;
    assign _418 = ~ _411;
    assign read_enable_14 = _102 & _418;
    assign write_enable_18 = _402 & _411;
    assign _420 = write_enable_18 | read_enable_14;
    assign address_19 = _411 ? _164 : _137;
    assign _413 = ~ _411;
    assign read_enable_15 = _102 & _413;
    assign _411 = ~ PHASE_3;
    assign write_enable_19 = _395 & _411;
    assign _415 = write_enable_19 | read_enable_15;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_8
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_415), .regcea(vdd), .wea(write_enable_19), .addra(address_19), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_420), .regceb(vdd), .web(write_enable_18), .addrb(address_18), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_423[131:131]), .sbiterrb(_423[130:130]), .doutb(_423[129:66]), .dbiterra(_423[65:65]), .sbiterra(_423[64:64]), .douta(_423[63:0]) );
    assign _424 = _423[63:0];
    assign _491 = _490[127:64];
    assign data_15 = _491;
    assign address_20 = PHASE_3 ? _199 : _172;
    assign _404 = ~ PHASE_3;
    assign read_enable_16 = _102 & _404;
    assign _401 = ~ _130;
    assign _402 = _129 & _401;
    assign write_enable_20 = _402 & PHASE_3;
    assign _406 = write_enable_20 | read_enable_16;
    assign address_21 = PHASE_3 ? _164 : _137;
    assign _397 = ~ PHASE_3;
    assign read_enable_17 = _102 & _397;
    assign _394 = ~ _130;
    assign _395 = _129 & _394;
    assign write_enable_21 = _395 & PHASE_3;
    assign _399 = write_enable_21 | read_enable_17;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_9
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_399), .regcea(vdd), .wea(write_enable_21), .addra(address_21), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_406), .regceb(vdd), .web(write_enable_20), .addrb(address_20), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_409[131:131]), .sbiterrb(_409[130:130]), .doutb(_409[129:66]), .dbiterra(_409[65:65]), .sbiterra(_409[64:64]), .douta(_409[63:0]) );
    assign _410 = _409[63:0];
    assign _492 = ~ PHASE_3;
    assign _13 = _492;
    always @(posedge _84) begin
        if (_82)
            PHASE_3 <= _392;
        else
            if (_99)
                PHASE_3 <= _13;
    end
    assign q0_0 = PHASE_3 ? _424 : _410;
    always @(posedge _84) begin
        if (_82)
            _390 <= _389;
        else
            _390 <= _92;
    end
    assign _481 = _390 ? _480 : q0_0;
    dp_29
        dp_5
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_481), .d2(_488), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_490[191:128]), .q2(_490[127:64]), .q1(_490[63:0]) );
    assign _493 = _490[63:0];
    assign data_19 = _493;
    assign address_22 = PHASE_4 ? _164 : _68;
    assign _557 = ~ PHASE_4;
    assign _556 = _70[6:6];
    assign read_enable_18 = _556 & _557;
    always @(posedge _84) begin
        if (_82)
            _527 <= _526;
        else
            _527 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _530 <= _529;
        else
            _530 <= _527;
    end
    always @(posedge _84) begin
        if (_82)
            _533 <= _532;
        else
            _533 <= _530;
    end
    always @(posedge _84) begin
        if (_82)
            _536 <= _535;
        else
            _536 <= _533;
    end
    always @(posedge _84) begin
        if (_82)
            _539 <= _538;
        else
            _539 <= _536;
    end
    always @(posedge _84) begin
        if (_82)
            _542 <= _541;
        else
            _542 <= _539;
    end
    always @(posedge _84) begin
        if (_82)
            _545 <= _544;
        else
            _545 <= _542;
    end
    always @(posedge _84) begin
        if (_82)
            _548 <= _547;
        else
            _548 <= _545;
    end
    always @(posedge _84) begin
        if (_82)
            _551 <= _550;
        else
            _551 <= _548;
    end
    assign _552 = ~ _551;
    always @(posedge _84) begin
        if (_82)
            _500 <= _499;
        else
            _500 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _503 <= _502;
        else
            _503 <= _500;
    end
    always @(posedge _84) begin
        if (_82)
            _506 <= _505;
        else
            _506 <= _503;
    end
    always @(posedge _84) begin
        if (_82)
            _509 <= _508;
        else
            _509 <= _506;
    end
    always @(posedge _84) begin
        if (_82)
            _512 <= _511;
        else
            _512 <= _509;
    end
    always @(posedge _84) begin
        if (_82)
            _515 <= _514;
        else
            _515 <= _512;
    end
    always @(posedge _84) begin
        if (_82)
            _518 <= _517;
        else
            _518 <= _515;
    end
    always @(posedge _84) begin
        if (_82)
            _521 <= _520;
        else
            _521 <= _518;
    end
    always @(posedge _84) begin
        if (_82)
            _524 <= _523;
        else
            _524 <= _521;
    end
    assign _553 = _524 & _552;
    assign _554 = _129 & _553;
    assign write_enable_22 = _554 & PHASE_4;
    assign _559 = write_enable_22 | read_enable_18;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_10
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_559), .regcea(vdd), .wea(write_enable_22), .addra(address_22), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_13), .regceb(vdd), .web(write_enable_13), .addrb(address_13), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_566[131:131]), .sbiterrb(_566[130:130]), .doutb(_566[129:66]), .dbiterra(_566[65:65]), .sbiterra(_566[64:64]), .douta(_566[63:0]) );
    assign _567 = _566[63:0];
    assign _497 = ~ PHASE_4;
    assign _15 = _497;
    always @(posedge _84) begin
        if (_82)
            PHASE_4 <= _495;
        else
            if (_72)
                PHASE_4 <= _15;
    end
    assign _579 = PHASE_4 ? _578 : _567;
    assign address_23 = _764 ? _199 : _759;
    assign write_enable_23 = _757 & _764;
    assign address_24 = _764 ? _164 : _68;
    assign _766 = ~ _764;
    assign read_enable_19 = _752 & _766;
    assign _764 = ~ PHASE_7;
    assign write_enable_24 = _750 & _764;
    assign _768 = write_enable_24 | read_enable_19;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_11
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_768), .regcea(vdd), .wea(write_enable_24), .addra(address_24), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_23), .regceb(vdd), .web(write_enable_23), .addrb(address_23), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_773[131:131]), .sbiterrb(_773[130:130]), .doutb(_773[129:66]), .dbiterra(_773[65:65]), .sbiterra(_773[64:64]), .douta(_773[63:0]) );
    assign _774 = _773[63:0];
    assign address_25 = PHASE_7 ? _199 : _759;
    assign _757 = _129 & _720;
    assign write_enable_25 = _757 & PHASE_7;
    assign _682 = _674[129:66];
    assign _681 = _661[129:66];
    assign _683 = PHASE_5 ? _682 : _681;
    assign _679 = _619[129:66];
    assign _678 = _605[129:66];
    assign q1_1 = PHASE_6 ? _679 : _678;
    assign _684 = _586 ? _683 : q1_1;
    assign address_26 = _663 ? _657 : _656;
    assign _669 = ~ _663;
    assign read_enable_20 = _102 & _669;
    assign address_27 = _663 ? _60 : _639;
    assign _665 = ~ _663;
    assign read_enable_21 = _102 & _665;
    assign _663 = ~ PHASE_5;
    assign write_enable_27 = _622 & _663;
    assign _667 = write_enable_27 | read_enable_21;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_12
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_667), .regcea(vdd), .wea(write_enable_27), .addra(address_27), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_20), .regceb(vdd), .web(write_enable_26), .addrb(address_26), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_674[131:131]), .sbiterrb(_674[130:130]), .doutb(_674[129:66]), .dbiterra(_674[65:65]), .sbiterra(_674[64:64]), .douta(_674[63:0]) );
    assign _675 = _674[63:0];
    assign _655 = _172[11:11];
    assign _654 = _172[10:10];
    assign _653 = _172[9:9];
    assign _652 = _172[8:8];
    assign _651 = _172[7:7];
    assign _650 = _172[6:6];
    assign _649 = _172[5:5];
    assign _648 = _172[4:4];
    assign _647 = _172[3:3];
    assign _646 = _172[2:2];
    assign _645 = _172[1:1];
    assign _644 = _172[0:0];
    assign _656 = { _644, _645, _646, _647, _648, _649, _650, _651, _652, _653, _654, _655 };
    assign address_28 = PHASE_5 ? _657 : _656;
    assign _641 = ~ PHASE_5;
    assign read_enable_22 = _102 & _641;
    assign data_25 = wr_d5;
    assign _638 = _137[11:11];
    assign _637 = _137[10:10];
    assign _636 = _137[9:9];
    assign _635 = _137[8:8];
    assign _634 = _137[7:7];
    assign _633 = _137[6:6];
    assign _632 = _137[5:5];
    assign _631 = _137[4:4];
    assign _630 = _137[3:3];
    assign _629 = _137[2:2];
    assign _628 = _137[1:1];
    assign _627 = _137[0:0];
    assign _639 = { _627, _628, _629, _630, _631, _632, _633, _634, _635, _636, _637, _638 };
    assign address_29 = PHASE_5 ? _60 : _639;
    assign _624 = ~ PHASE_5;
    assign read_enable_23 = _102 & _624;
    assign _622 = _62[5:5];
    assign write_enable_29 = _622 & PHASE_5;
    assign _626 = write_enable_29 | read_enable_23;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_13
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_626), .regcea(vdd), .wea(write_enable_29), .addra(address_29), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_22), .regceb(vdd), .web(write_enable_28), .addrb(address_28), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_661[131:131]), .sbiterrb(_661[130:130]), .doutb(_661[129:66]), .dbiterra(_661[65:65]), .sbiterra(_661[64:64]), .douta(_661[63:0]) );
    assign _662 = _661[63:0];
    assign _583 = ~ PHASE_5;
    assign _19 = _583;
    always @(posedge _84) begin
        if (_82)
            PHASE_5 <= _581;
        else
            if (_72)
                PHASE_5 <= _19;
    end
    assign _676 = PHASE_5 ? _675 : _662;
    assign address_30 = _607 ? _199 : _172;
    assign _614 = ~ _607;
    assign read_enable_24 = _102 & _614;
    assign write_enable_30 = _598 & _607;
    assign _616 = write_enable_30 | read_enable_24;
    assign address_31 = _607 ? _164 : _137;
    assign _609 = ~ _607;
    assign read_enable_25 = _102 & _609;
    assign _607 = ~ PHASE_6;
    assign write_enable_31 = _591 & _607;
    assign _611 = write_enable_31 | read_enable_25;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_14
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_611), .regcea(vdd), .wea(write_enable_31), .addra(address_31), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_616), .regceb(vdd), .web(write_enable_30), .addrb(address_30), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_619[131:131]), .sbiterrb(_619[130:130]), .doutb(_619[129:66]), .dbiterra(_619[65:65]), .sbiterra(_619[64:64]), .douta(_619[63:0]) );
    assign _620 = _619[63:0];
    assign _687 = _686[127:64];
    assign data_27 = _687;
    assign address_32 = PHASE_6 ? _199 : _172;
    assign _600 = ~ PHASE_6;
    assign read_enable_26 = _102 & _600;
    assign _597 = ~ _130;
    assign _598 = _129 & _597;
    assign write_enable_32 = _598 & PHASE_6;
    assign _602 = write_enable_32 | read_enable_26;
    assign address_33 = PHASE_6 ? _164 : _137;
    assign _593 = ~ PHASE_6;
    assign read_enable_27 = _102 & _593;
    assign _590 = ~ _130;
    assign _591 = _129 & _590;
    assign write_enable_33 = _591 & PHASE_6;
    assign _595 = write_enable_33 | read_enable_27;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_15
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_595), .regcea(vdd), .wea(write_enable_33), .addra(address_33), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_602), .regceb(vdd), .web(write_enable_32), .addrb(address_32), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_605[131:131]), .sbiterrb(_605[130:130]), .doutb(_605[129:66]), .dbiterra(_605[65:65]), .sbiterra(_605[64:64]), .douta(_605[63:0]) );
    assign _606 = _605[63:0];
    assign _688 = ~ PHASE_6;
    assign _21 = _688;
    always @(posedge _84) begin
        if (_82)
            PHASE_6 <= _588;
        else
            if (_99)
                PHASE_6 <= _21;
    end
    assign q0_1 = PHASE_6 ? _620 : _606;
    always @(posedge _84) begin
        if (_82)
            _586 <= _585;
        else
            _586 <= _92;
    end
    assign _677 = _586 ? _676 : q0_1;
    dp_28
        dp_4
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_677), .d2(_684), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_686[191:128]), .q2(_686[127:64]), .q1(_686[63:0]) );
    assign _689 = _686[63:0];
    assign data_31 = _689;
    assign address_34 = PHASE_7 ? _164 : _68;
    assign _753 = ~ PHASE_7;
    assign _752 = _70[5:5];
    assign read_enable_28 = _752 & _753;
    always @(posedge _84) begin
        if (_82)
            _723 <= _722;
        else
            _723 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _726 <= _725;
        else
            _726 <= _723;
    end
    always @(posedge _84) begin
        if (_82)
            _729 <= _728;
        else
            _729 <= _726;
    end
    always @(posedge _84) begin
        if (_82)
            _732 <= _731;
        else
            _732 <= _729;
    end
    always @(posedge _84) begin
        if (_82)
            _735 <= _734;
        else
            _735 <= _732;
    end
    always @(posedge _84) begin
        if (_82)
            _738 <= _737;
        else
            _738 <= _735;
    end
    always @(posedge _84) begin
        if (_82)
            _741 <= _740;
        else
            _741 <= _738;
    end
    always @(posedge _84) begin
        if (_82)
            _744 <= _743;
        else
            _744 <= _741;
    end
    always @(posedge _84) begin
        if (_82)
            _747 <= _746;
        else
            _747 <= _744;
    end
    assign _748 = ~ _747;
    always @(posedge _84) begin
        if (_82)
            _696 <= _695;
        else
            _696 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _699 <= _698;
        else
            _699 <= _696;
    end
    always @(posedge _84) begin
        if (_82)
            _702 <= _701;
        else
            _702 <= _699;
    end
    always @(posedge _84) begin
        if (_82)
            _705 <= _704;
        else
            _705 <= _702;
    end
    always @(posedge _84) begin
        if (_82)
            _708 <= _707;
        else
            _708 <= _705;
    end
    always @(posedge _84) begin
        if (_82)
            _711 <= _710;
        else
            _711 <= _708;
    end
    always @(posedge _84) begin
        if (_82)
            _714 <= _713;
        else
            _714 <= _711;
    end
    always @(posedge _84) begin
        if (_82)
            _717 <= _716;
        else
            _717 <= _714;
    end
    always @(posedge _84) begin
        if (_82)
            _720 <= _719;
        else
            _720 <= _717;
    end
    assign _749 = _720 & _748;
    assign _750 = _129 & _749;
    assign write_enable_34 = _750 & PHASE_7;
    assign _755 = write_enable_34 | read_enable_28;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_16
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_755), .regcea(vdd), .wea(write_enable_34), .addra(address_34), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_25), .regceb(vdd), .web(write_enable_25), .addrb(address_25), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_762[131:131]), .sbiterrb(_762[130:130]), .doutb(_762[129:66]), .dbiterra(_762[65:65]), .sbiterra(_762[64:64]), .douta(_762[63:0]) );
    assign _763 = _762[63:0];
    assign _693 = ~ PHASE_7;
    assign _23 = _693;
    always @(posedge _84) begin
        if (_82)
            PHASE_7 <= _691;
        else
            if (_72)
                PHASE_7 <= _23;
    end
    assign _775 = PHASE_7 ? _774 : _763;
    assign address_35 = _960 ? _199 : _955;
    assign write_enable_35 = _953 & _960;
    assign address_36 = _960 ? _164 : _68;
    assign _962 = ~ _960;
    assign read_enable_29 = _948 & _962;
    assign _960 = ~ PHASE_10;
    assign write_enable_36 = _946 & _960;
    assign _964 = write_enable_36 | read_enable_29;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_17
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_964), .regcea(vdd), .wea(write_enable_36), .addra(address_36), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_35), .regceb(vdd), .web(write_enable_35), .addrb(address_35), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_969[131:131]), .sbiterrb(_969[130:130]), .doutb(_969[129:66]), .dbiterra(_969[65:65]), .sbiterra(_969[64:64]), .douta(_969[63:0]) );
    assign _970 = _969[63:0];
    assign address_37 = PHASE_10 ? _199 : _955;
    assign _953 = _129 & _916;
    assign write_enable_37 = _953 & PHASE_10;
    assign _878 = _870[129:66];
    assign _877 = _857[129:66];
    assign _879 = PHASE_8 ? _878 : _877;
    assign _875 = _815[129:66];
    assign _874 = _801[129:66];
    assign q1_2 = PHASE_9 ? _875 : _874;
    assign _880 = _782 ? _879 : q1_2;
    assign address_38 = _859 ? _853 : _852;
    assign _865 = ~ _859;
    assign read_enable_30 = _102 & _865;
    assign address_39 = _859 ? _60 : _835;
    assign _861 = ~ _859;
    assign read_enable_31 = _102 & _861;
    assign _859 = ~ PHASE_8;
    assign write_enable_39 = _818 & _859;
    assign _863 = write_enable_39 | read_enable_31;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_18
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_863), .regcea(vdd), .wea(write_enable_39), .addra(address_39), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_30), .regceb(vdd), .web(write_enable_38), .addrb(address_38), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_870[131:131]), .sbiterrb(_870[130:130]), .doutb(_870[129:66]), .dbiterra(_870[65:65]), .sbiterra(_870[64:64]), .douta(_870[63:0]) );
    assign _871 = _870[63:0];
    assign _851 = _172[11:11];
    assign _850 = _172[10:10];
    assign _849 = _172[9:9];
    assign _848 = _172[8:8];
    assign _847 = _172[7:7];
    assign _846 = _172[6:6];
    assign _845 = _172[5:5];
    assign _844 = _172[4:4];
    assign _843 = _172[3:3];
    assign _842 = _172[2:2];
    assign _841 = _172[1:1];
    assign _840 = _172[0:0];
    assign _852 = { _840, _841, _842, _843, _844, _845, _846, _847, _848, _849, _850, _851 };
    assign address_40 = PHASE_8 ? _853 : _852;
    assign _837 = ~ PHASE_8;
    assign read_enable_32 = _102 & _837;
    assign data_37 = wr_d4;
    assign _834 = _137[11:11];
    assign _833 = _137[10:10];
    assign _832 = _137[9:9];
    assign _831 = _137[8:8];
    assign _830 = _137[7:7];
    assign _829 = _137[6:6];
    assign _828 = _137[5:5];
    assign _827 = _137[4:4];
    assign _826 = _137[3:3];
    assign _825 = _137[2:2];
    assign _824 = _137[1:1];
    assign _823 = _137[0:0];
    assign _835 = { _823, _824, _825, _826, _827, _828, _829, _830, _831, _832, _833, _834 };
    assign address_41 = PHASE_8 ? _60 : _835;
    assign _820 = ~ PHASE_8;
    assign read_enable_33 = _102 & _820;
    assign _818 = _62[4:4];
    assign write_enable_41 = _818 & PHASE_8;
    assign _822 = write_enable_41 | read_enable_33;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_19
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_822), .regcea(vdd), .wea(write_enable_41), .addra(address_41), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_32), .regceb(vdd), .web(write_enable_40), .addrb(address_40), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_857[131:131]), .sbiterrb(_857[130:130]), .doutb(_857[129:66]), .dbiterra(_857[65:65]), .sbiterra(_857[64:64]), .douta(_857[63:0]) );
    assign _858 = _857[63:0];
    assign _779 = ~ PHASE_8;
    assign _27 = _779;
    always @(posedge _84) begin
        if (_82)
            PHASE_8 <= _777;
        else
            if (_72)
                PHASE_8 <= _27;
    end
    assign _872 = PHASE_8 ? _871 : _858;
    assign address_42 = _803 ? _199 : _172;
    assign _810 = ~ _803;
    assign read_enable_34 = _102 & _810;
    assign write_enable_42 = _794 & _803;
    assign _812 = write_enable_42 | read_enable_34;
    assign address_43 = _803 ? _164 : _137;
    assign _805 = ~ _803;
    assign read_enable_35 = _102 & _805;
    assign _803 = ~ PHASE_9;
    assign write_enable_43 = _787 & _803;
    assign _807 = write_enable_43 | read_enable_35;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_20
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_807), .regcea(vdd), .wea(write_enable_43), .addra(address_43), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_812), .regceb(vdd), .web(write_enable_42), .addrb(address_42), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_815[131:131]), .sbiterrb(_815[130:130]), .doutb(_815[129:66]), .dbiterra(_815[65:65]), .sbiterra(_815[64:64]), .douta(_815[63:0]) );
    assign _816 = _815[63:0];
    assign _883 = _882[127:64];
    assign data_39 = _883;
    assign address_44 = PHASE_9 ? _199 : _172;
    assign _796 = ~ PHASE_9;
    assign read_enable_36 = _102 & _796;
    assign _793 = ~ _130;
    assign _794 = _129 & _793;
    assign write_enable_44 = _794 & PHASE_9;
    assign _798 = write_enable_44 | read_enable_36;
    assign address_45 = PHASE_9 ? _164 : _137;
    assign _789 = ~ PHASE_9;
    assign read_enable_37 = _102 & _789;
    assign _786 = ~ _130;
    assign _787 = _129 & _786;
    assign write_enable_45 = _787 & PHASE_9;
    assign _791 = write_enable_45 | read_enable_37;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_21
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_791), .regcea(vdd), .wea(write_enable_45), .addra(address_45), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_798), .regceb(vdd), .web(write_enable_44), .addrb(address_44), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_801[131:131]), .sbiterrb(_801[130:130]), .doutb(_801[129:66]), .dbiterra(_801[65:65]), .sbiterra(_801[64:64]), .douta(_801[63:0]) );
    assign _802 = _801[63:0];
    assign _884 = ~ PHASE_9;
    assign _29 = _884;
    always @(posedge _84) begin
        if (_82)
            PHASE_9 <= _784;
        else
            if (_99)
                PHASE_9 <= _29;
    end
    assign q0_2 = PHASE_9 ? _816 : _802;
    always @(posedge _84) begin
        if (_82)
            _782 <= _781;
        else
            _782 <= _92;
    end
    assign _873 = _782 ? _872 : q0_2;
    dp_27
        dp_3
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_873), .d2(_880), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_882[191:128]), .q2(_882[127:64]), .q1(_882[63:0]) );
    assign _885 = _882[63:0];
    assign data_43 = _885;
    assign address_46 = PHASE_10 ? _164 : _68;
    assign _949 = ~ PHASE_10;
    assign _948 = _70[4:4];
    assign read_enable_38 = _948 & _949;
    always @(posedge _84) begin
        if (_82)
            _919 <= _918;
        else
            _919 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _922 <= _921;
        else
            _922 <= _919;
    end
    always @(posedge _84) begin
        if (_82)
            _925 <= _924;
        else
            _925 <= _922;
    end
    always @(posedge _84) begin
        if (_82)
            _928 <= _927;
        else
            _928 <= _925;
    end
    always @(posedge _84) begin
        if (_82)
            _931 <= _930;
        else
            _931 <= _928;
    end
    always @(posedge _84) begin
        if (_82)
            _934 <= _933;
        else
            _934 <= _931;
    end
    always @(posedge _84) begin
        if (_82)
            _937 <= _936;
        else
            _937 <= _934;
    end
    always @(posedge _84) begin
        if (_82)
            _940 <= _939;
        else
            _940 <= _937;
    end
    always @(posedge _84) begin
        if (_82)
            _943 <= _942;
        else
            _943 <= _940;
    end
    assign _944 = ~ _943;
    always @(posedge _84) begin
        if (_82)
            _892 <= _891;
        else
            _892 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _895 <= _894;
        else
            _895 <= _892;
    end
    always @(posedge _84) begin
        if (_82)
            _898 <= _897;
        else
            _898 <= _895;
    end
    always @(posedge _84) begin
        if (_82)
            _901 <= _900;
        else
            _901 <= _898;
    end
    always @(posedge _84) begin
        if (_82)
            _904 <= _903;
        else
            _904 <= _901;
    end
    always @(posedge _84) begin
        if (_82)
            _907 <= _906;
        else
            _907 <= _904;
    end
    always @(posedge _84) begin
        if (_82)
            _910 <= _909;
        else
            _910 <= _907;
    end
    always @(posedge _84) begin
        if (_82)
            _913 <= _912;
        else
            _913 <= _910;
    end
    always @(posedge _84) begin
        if (_82)
            _916 <= _915;
        else
            _916 <= _913;
    end
    assign _945 = _916 & _944;
    assign _946 = _129 & _945;
    assign write_enable_46 = _946 & PHASE_10;
    assign _951 = write_enable_46 | read_enable_38;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_22
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_951), .regcea(vdd), .wea(write_enable_46), .addra(address_46), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_37), .regceb(vdd), .web(write_enable_37), .addrb(address_37), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_958[131:131]), .sbiterrb(_958[130:130]), .doutb(_958[129:66]), .dbiterra(_958[65:65]), .sbiterra(_958[64:64]), .douta(_958[63:0]) );
    assign _959 = _958[63:0];
    assign _889 = ~ PHASE_10;
    assign _31 = _889;
    always @(posedge _84) begin
        if (_82)
            PHASE_10 <= _887;
        else
            if (_72)
                PHASE_10 <= _31;
    end
    assign _971 = PHASE_10 ? _970 : _959;
    assign address_47 = _1156 ? _199 : _1151;
    assign write_enable_47 = _1149 & _1156;
    assign address_48 = _1156 ? _164 : _68;
    assign _1158 = ~ _1156;
    assign read_enable_39 = _1144 & _1158;
    assign _1156 = ~ PHASE_13;
    assign write_enable_48 = _1142 & _1156;
    assign _1160 = write_enable_48 | read_enable_39;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_23
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1160), .regcea(vdd), .wea(write_enable_48), .addra(address_48), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_47), .regceb(vdd), .web(write_enable_47), .addrb(address_47), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1165[131:131]), .sbiterrb(_1165[130:130]), .doutb(_1165[129:66]), .dbiterra(_1165[65:65]), .sbiterra(_1165[64:64]), .douta(_1165[63:0]) );
    assign _1166 = _1165[63:0];
    assign address_49 = PHASE_13 ? _199 : _1151;
    assign _1149 = _129 & _1112;
    assign write_enable_49 = _1149 & PHASE_13;
    assign _1074 = _1066[129:66];
    assign _1073 = _1053[129:66];
    assign _1075 = PHASE_11 ? _1074 : _1073;
    assign _1071 = _1011[129:66];
    assign _1070 = _997[129:66];
    assign q1_3 = PHASE_12 ? _1071 : _1070;
    assign _1076 = _978 ? _1075 : q1_3;
    assign address_50 = _1055 ? _1049 : _1048;
    assign _1061 = ~ _1055;
    assign read_enable_40 = _102 & _1061;
    assign address_51 = _1055 ? _60 : _1031;
    assign _1057 = ~ _1055;
    assign read_enable_41 = _102 & _1057;
    assign _1055 = ~ PHASE_11;
    assign write_enable_51 = _1014 & _1055;
    assign _1059 = write_enable_51 | read_enable_41;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_24
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1059), .regcea(vdd), .wea(write_enable_51), .addra(address_51), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_40), .regceb(vdd), .web(write_enable_50), .addrb(address_50), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1066[131:131]), .sbiterrb(_1066[130:130]), .doutb(_1066[129:66]), .dbiterra(_1066[65:65]), .sbiterra(_1066[64:64]), .douta(_1066[63:0]) );
    assign _1067 = _1066[63:0];
    assign _1047 = _172[11:11];
    assign _1046 = _172[10:10];
    assign _1045 = _172[9:9];
    assign _1044 = _172[8:8];
    assign _1043 = _172[7:7];
    assign _1042 = _172[6:6];
    assign _1041 = _172[5:5];
    assign _1040 = _172[4:4];
    assign _1039 = _172[3:3];
    assign _1038 = _172[2:2];
    assign _1037 = _172[1:1];
    assign _1036 = _172[0:0];
    assign _1048 = { _1036, _1037, _1038, _1039, _1040, _1041, _1042, _1043, _1044, _1045, _1046, _1047 };
    assign address_52 = PHASE_11 ? _1049 : _1048;
    assign _1033 = ~ PHASE_11;
    assign read_enable_42 = _102 & _1033;
    assign data_49 = wr_d3;
    assign _1030 = _137[11:11];
    assign _1029 = _137[10:10];
    assign _1028 = _137[9:9];
    assign _1027 = _137[8:8];
    assign _1026 = _137[7:7];
    assign _1025 = _137[6:6];
    assign _1024 = _137[5:5];
    assign _1023 = _137[4:4];
    assign _1022 = _137[3:3];
    assign _1021 = _137[2:2];
    assign _1020 = _137[1:1];
    assign _1019 = _137[0:0];
    assign _1031 = { _1019, _1020, _1021, _1022, _1023, _1024, _1025, _1026, _1027, _1028, _1029, _1030 };
    assign address_53 = PHASE_11 ? _60 : _1031;
    assign _1016 = ~ PHASE_11;
    assign read_enable_43 = _102 & _1016;
    assign _1014 = _62[3:3];
    assign write_enable_53 = _1014 & PHASE_11;
    assign _1018 = write_enable_53 | read_enable_43;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_25
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1018), .regcea(vdd), .wea(write_enable_53), .addra(address_53), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_42), .regceb(vdd), .web(write_enable_52), .addrb(address_52), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1053[131:131]), .sbiterrb(_1053[130:130]), .doutb(_1053[129:66]), .dbiterra(_1053[65:65]), .sbiterra(_1053[64:64]), .douta(_1053[63:0]) );
    assign _1054 = _1053[63:0];
    assign _975 = ~ PHASE_11;
    assign _35 = _975;
    always @(posedge _84) begin
        if (_82)
            PHASE_11 <= _973;
        else
            if (_72)
                PHASE_11 <= _35;
    end
    assign _1068 = PHASE_11 ? _1067 : _1054;
    assign address_54 = _999 ? _199 : _172;
    assign _1006 = ~ _999;
    assign read_enable_44 = _102 & _1006;
    assign write_enable_54 = _990 & _999;
    assign _1008 = write_enable_54 | read_enable_44;
    assign address_55 = _999 ? _164 : _137;
    assign _1001 = ~ _999;
    assign read_enable_45 = _102 & _1001;
    assign _999 = ~ PHASE_12;
    assign write_enable_55 = _983 & _999;
    assign _1003 = write_enable_55 | read_enable_45;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_26
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1003), .regcea(vdd), .wea(write_enable_55), .addra(address_55), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1008), .regceb(vdd), .web(write_enable_54), .addrb(address_54), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1011[131:131]), .sbiterrb(_1011[130:130]), .doutb(_1011[129:66]), .dbiterra(_1011[65:65]), .sbiterra(_1011[64:64]), .douta(_1011[63:0]) );
    assign _1012 = _1011[63:0];
    assign _1079 = _1078[127:64];
    assign data_51 = _1079;
    assign address_56 = PHASE_12 ? _199 : _172;
    assign _992 = ~ PHASE_12;
    assign read_enable_46 = _102 & _992;
    assign _989 = ~ _130;
    assign _990 = _129 & _989;
    assign write_enable_56 = _990 & PHASE_12;
    assign _994 = write_enable_56 | read_enable_46;
    assign address_57 = PHASE_12 ? _164 : _137;
    assign _985 = ~ PHASE_12;
    assign read_enable_47 = _102 & _985;
    assign _982 = ~ _130;
    assign _983 = _129 & _982;
    assign write_enable_57 = _983 & PHASE_12;
    assign _987 = write_enable_57 | read_enable_47;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_27
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_987), .regcea(vdd), .wea(write_enable_57), .addra(address_57), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_994), .regceb(vdd), .web(write_enable_56), .addrb(address_56), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_997[131:131]), .sbiterrb(_997[130:130]), .doutb(_997[129:66]), .dbiterra(_997[65:65]), .sbiterra(_997[64:64]), .douta(_997[63:0]) );
    assign _998 = _997[63:0];
    assign _1080 = ~ PHASE_12;
    assign _37 = _1080;
    always @(posedge _84) begin
        if (_82)
            PHASE_12 <= _980;
        else
            if (_99)
                PHASE_12 <= _37;
    end
    assign q0_3 = PHASE_12 ? _1012 : _998;
    always @(posedge _84) begin
        if (_82)
            _978 <= _977;
        else
            _978 <= _92;
    end
    assign _1069 = _978 ? _1068 : q0_3;
    dp_26
        dp_2
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1069), .d2(_1076), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1078[191:128]), .q2(_1078[127:64]), .q1(_1078[63:0]) );
    assign _1081 = _1078[63:0];
    assign data_55 = _1081;
    assign address_58 = PHASE_13 ? _164 : _68;
    assign _1145 = ~ PHASE_13;
    assign _1144 = _70[3:3];
    assign read_enable_48 = _1144 & _1145;
    always @(posedge _84) begin
        if (_82)
            _1115 <= _1114;
        else
            _1115 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1118 <= _1117;
        else
            _1118 <= _1115;
    end
    always @(posedge _84) begin
        if (_82)
            _1121 <= _1120;
        else
            _1121 <= _1118;
    end
    always @(posedge _84) begin
        if (_82)
            _1124 <= _1123;
        else
            _1124 <= _1121;
    end
    always @(posedge _84) begin
        if (_82)
            _1127 <= _1126;
        else
            _1127 <= _1124;
    end
    always @(posedge _84) begin
        if (_82)
            _1130 <= _1129;
        else
            _1130 <= _1127;
    end
    always @(posedge _84) begin
        if (_82)
            _1133 <= _1132;
        else
            _1133 <= _1130;
    end
    always @(posedge _84) begin
        if (_82)
            _1136 <= _1135;
        else
            _1136 <= _1133;
    end
    always @(posedge _84) begin
        if (_82)
            _1139 <= _1138;
        else
            _1139 <= _1136;
    end
    assign _1140 = ~ _1139;
    always @(posedge _84) begin
        if (_82)
            _1088 <= _1087;
        else
            _1088 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1091 <= _1090;
        else
            _1091 <= _1088;
    end
    always @(posedge _84) begin
        if (_82)
            _1094 <= _1093;
        else
            _1094 <= _1091;
    end
    always @(posedge _84) begin
        if (_82)
            _1097 <= _1096;
        else
            _1097 <= _1094;
    end
    always @(posedge _84) begin
        if (_82)
            _1100 <= _1099;
        else
            _1100 <= _1097;
    end
    always @(posedge _84) begin
        if (_82)
            _1103 <= _1102;
        else
            _1103 <= _1100;
    end
    always @(posedge _84) begin
        if (_82)
            _1106 <= _1105;
        else
            _1106 <= _1103;
    end
    always @(posedge _84) begin
        if (_82)
            _1109 <= _1108;
        else
            _1109 <= _1106;
    end
    always @(posedge _84) begin
        if (_82)
            _1112 <= _1111;
        else
            _1112 <= _1109;
    end
    assign _1141 = _1112 & _1140;
    assign _1142 = _129 & _1141;
    assign write_enable_58 = _1142 & PHASE_13;
    assign _1147 = write_enable_58 | read_enable_48;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_28
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1147), .regcea(vdd), .wea(write_enable_58), .addra(address_58), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_49), .regceb(vdd), .web(write_enable_49), .addrb(address_49), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1154[131:131]), .sbiterrb(_1154[130:130]), .doutb(_1154[129:66]), .dbiterra(_1154[65:65]), .sbiterra(_1154[64:64]), .douta(_1154[63:0]) );
    assign _1155 = _1154[63:0];
    assign _1085 = ~ PHASE_13;
    assign _39 = _1085;
    always @(posedge _84) begin
        if (_82)
            PHASE_13 <= _1083;
        else
            if (_72)
                PHASE_13 <= _39;
    end
    assign _1167 = PHASE_13 ? _1166 : _1155;
    assign address_59 = _1352 ? _199 : _1347;
    assign write_enable_59 = _1345 & _1352;
    assign address_60 = _1352 ? _164 : _68;
    assign _1354 = ~ _1352;
    assign read_enable_49 = _1340 & _1354;
    assign _1352 = ~ PHASE_16;
    assign write_enable_60 = _1338 & _1352;
    assign _1356 = write_enable_60 | read_enable_49;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_29
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1356), .regcea(vdd), .wea(write_enable_60), .addra(address_60), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_59), .regceb(vdd), .web(write_enable_59), .addrb(address_59), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1361[131:131]), .sbiterrb(_1361[130:130]), .doutb(_1361[129:66]), .dbiterra(_1361[65:65]), .sbiterra(_1361[64:64]), .douta(_1361[63:0]) );
    assign _1362 = _1361[63:0];
    assign address_61 = PHASE_16 ? _199 : _1347;
    assign _1345 = _129 & _1308;
    assign write_enable_61 = _1345 & PHASE_16;
    assign _1270 = _1262[129:66];
    assign _1269 = _1249[129:66];
    assign _1271 = PHASE_14 ? _1270 : _1269;
    assign _1267 = _1207[129:66];
    assign _1266 = _1193[129:66];
    assign q1_4 = PHASE_15 ? _1267 : _1266;
    assign _1272 = _1174 ? _1271 : q1_4;
    assign address_62 = _1251 ? _1245 : _1244;
    assign _1257 = ~ _1251;
    assign read_enable_50 = _102 & _1257;
    assign address_63 = _1251 ? _60 : _1227;
    assign _1253 = ~ _1251;
    assign read_enable_51 = _102 & _1253;
    assign _1251 = ~ PHASE_14;
    assign write_enable_63 = _1210 & _1251;
    assign _1255 = write_enable_63 | read_enable_51;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_30
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1255), .regcea(vdd), .wea(write_enable_63), .addra(address_63), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_50), .regceb(vdd), .web(write_enable_62), .addrb(address_62), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1262[131:131]), .sbiterrb(_1262[130:130]), .doutb(_1262[129:66]), .dbiterra(_1262[65:65]), .sbiterra(_1262[64:64]), .douta(_1262[63:0]) );
    assign _1263 = _1262[63:0];
    assign _1243 = _172[11:11];
    assign _1242 = _172[10:10];
    assign _1241 = _172[9:9];
    assign _1240 = _172[8:8];
    assign _1239 = _172[7:7];
    assign _1238 = _172[6:6];
    assign _1237 = _172[5:5];
    assign _1236 = _172[4:4];
    assign _1235 = _172[3:3];
    assign _1234 = _172[2:2];
    assign _1233 = _172[1:1];
    assign _1232 = _172[0:0];
    assign _1244 = { _1232, _1233, _1234, _1235, _1236, _1237, _1238, _1239, _1240, _1241, _1242, _1243 };
    assign address_64 = PHASE_14 ? _1245 : _1244;
    assign _1229 = ~ PHASE_14;
    assign read_enable_52 = _102 & _1229;
    assign data_61 = wr_d2;
    assign _1226 = _137[11:11];
    assign _1225 = _137[10:10];
    assign _1224 = _137[9:9];
    assign _1223 = _137[8:8];
    assign _1222 = _137[7:7];
    assign _1221 = _137[6:6];
    assign _1220 = _137[5:5];
    assign _1219 = _137[4:4];
    assign _1218 = _137[3:3];
    assign _1217 = _137[2:2];
    assign _1216 = _137[1:1];
    assign _1215 = _137[0:0];
    assign _1227 = { _1215, _1216, _1217, _1218, _1219, _1220, _1221, _1222, _1223, _1224, _1225, _1226 };
    assign address_65 = PHASE_14 ? _60 : _1227;
    assign _1212 = ~ PHASE_14;
    assign read_enable_53 = _102 & _1212;
    assign _1210 = _62[2:2];
    assign write_enable_65 = _1210 & PHASE_14;
    assign _1214 = write_enable_65 | read_enable_53;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_31
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1214), .regcea(vdd), .wea(write_enable_65), .addra(address_65), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_52), .regceb(vdd), .web(write_enable_64), .addrb(address_64), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1249[131:131]), .sbiterrb(_1249[130:130]), .doutb(_1249[129:66]), .dbiterra(_1249[65:65]), .sbiterra(_1249[64:64]), .douta(_1249[63:0]) );
    assign _1250 = _1249[63:0];
    assign _1171 = ~ PHASE_14;
    assign _43 = _1171;
    always @(posedge _84) begin
        if (_82)
            PHASE_14 <= _1169;
        else
            if (_72)
                PHASE_14 <= _43;
    end
    assign _1264 = PHASE_14 ? _1263 : _1250;
    assign address_66 = _1195 ? _199 : _172;
    assign _1202 = ~ _1195;
    assign read_enable_54 = _102 & _1202;
    assign write_enable_66 = _1186 & _1195;
    assign _1204 = write_enable_66 | read_enable_54;
    assign address_67 = _1195 ? _164 : _137;
    assign _1197 = ~ _1195;
    assign read_enable_55 = _102 & _1197;
    assign _1195 = ~ PHASE_15;
    assign write_enable_67 = _1179 & _1195;
    assign _1199 = write_enable_67 | read_enable_55;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_32
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1199), .regcea(vdd), .wea(write_enable_67), .addra(address_67), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1204), .regceb(vdd), .web(write_enable_66), .addrb(address_66), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1207[131:131]), .sbiterrb(_1207[130:130]), .doutb(_1207[129:66]), .dbiterra(_1207[65:65]), .sbiterra(_1207[64:64]), .douta(_1207[63:0]) );
    assign _1208 = _1207[63:0];
    assign _1275 = _1274[127:64];
    assign data_63 = _1275;
    assign address_68 = PHASE_15 ? _199 : _172;
    assign _1188 = ~ PHASE_15;
    assign read_enable_56 = _102 & _1188;
    assign _1185 = ~ _130;
    assign _1186 = _129 & _1185;
    assign write_enable_68 = _1186 & PHASE_15;
    assign _1190 = write_enable_68 | read_enable_56;
    assign address_69 = PHASE_15 ? _164 : _137;
    assign _1181 = ~ PHASE_15;
    assign read_enable_57 = _102 & _1181;
    assign _1178 = ~ _130;
    assign _1179 = _129 & _1178;
    assign write_enable_69 = _1179 & PHASE_15;
    assign _1183 = write_enable_69 | read_enable_57;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_33
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1183), .regcea(vdd), .wea(write_enable_69), .addra(address_69), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1190), .regceb(vdd), .web(write_enable_68), .addrb(address_68), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1193[131:131]), .sbiterrb(_1193[130:130]), .doutb(_1193[129:66]), .dbiterra(_1193[65:65]), .sbiterra(_1193[64:64]), .douta(_1193[63:0]) );
    assign _1194 = _1193[63:0];
    assign _1276 = ~ PHASE_15;
    assign _45 = _1276;
    always @(posedge _84) begin
        if (_82)
            PHASE_15 <= _1176;
        else
            if (_99)
                PHASE_15 <= _45;
    end
    assign q0_4 = PHASE_15 ? _1208 : _1194;
    always @(posedge _84) begin
        if (_82)
            _1174 <= _1173;
        else
            _1174 <= _92;
    end
    assign _1265 = _1174 ? _1264 : q0_4;
    dp_25
        dp_1
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1265), .d2(_1272), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1274[191:128]), .q2(_1274[127:64]), .q1(_1274[63:0]) );
    assign _1277 = _1274[63:0];
    assign data_67 = _1277;
    assign address_70 = PHASE_16 ? _164 : _68;
    assign _1341 = ~ PHASE_16;
    assign _1340 = _70[2:2];
    assign read_enable_58 = _1340 & _1341;
    always @(posedge _84) begin
        if (_82)
            _1311 <= _1310;
        else
            _1311 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1314 <= _1313;
        else
            _1314 <= _1311;
    end
    always @(posedge _84) begin
        if (_82)
            _1317 <= _1316;
        else
            _1317 <= _1314;
    end
    always @(posedge _84) begin
        if (_82)
            _1320 <= _1319;
        else
            _1320 <= _1317;
    end
    always @(posedge _84) begin
        if (_82)
            _1323 <= _1322;
        else
            _1323 <= _1320;
    end
    always @(posedge _84) begin
        if (_82)
            _1326 <= _1325;
        else
            _1326 <= _1323;
    end
    always @(posedge _84) begin
        if (_82)
            _1329 <= _1328;
        else
            _1329 <= _1326;
    end
    always @(posedge _84) begin
        if (_82)
            _1332 <= _1331;
        else
            _1332 <= _1329;
    end
    always @(posedge _84) begin
        if (_82)
            _1335 <= _1334;
        else
            _1335 <= _1332;
    end
    assign _1336 = ~ _1335;
    always @(posedge _84) begin
        if (_82)
            _1284 <= _1283;
        else
            _1284 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1287 <= _1286;
        else
            _1287 <= _1284;
    end
    always @(posedge _84) begin
        if (_82)
            _1290 <= _1289;
        else
            _1290 <= _1287;
    end
    always @(posedge _84) begin
        if (_82)
            _1293 <= _1292;
        else
            _1293 <= _1290;
    end
    always @(posedge _84) begin
        if (_82)
            _1296 <= _1295;
        else
            _1296 <= _1293;
    end
    always @(posedge _84) begin
        if (_82)
            _1299 <= _1298;
        else
            _1299 <= _1296;
    end
    always @(posedge _84) begin
        if (_82)
            _1302 <= _1301;
        else
            _1302 <= _1299;
    end
    always @(posedge _84) begin
        if (_82)
            _1305 <= _1304;
        else
            _1305 <= _1302;
    end
    always @(posedge _84) begin
        if (_82)
            _1308 <= _1307;
        else
            _1308 <= _1305;
    end
    assign _1337 = _1308 & _1336;
    assign _1338 = _129 & _1337;
    assign write_enable_70 = _1338 & PHASE_16;
    assign _1343 = write_enable_70 | read_enable_58;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_34
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1343), .regcea(vdd), .wea(write_enable_70), .addra(address_70), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_61), .regceb(vdd), .web(write_enable_61), .addrb(address_61), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1350[131:131]), .sbiterrb(_1350[130:130]), .doutb(_1350[129:66]), .dbiterra(_1350[65:65]), .sbiterra(_1350[64:64]), .douta(_1350[63:0]) );
    assign _1351 = _1350[63:0];
    assign _1281 = ~ PHASE_16;
    assign _47 = _1281;
    always @(posedge _84) begin
        if (_82)
            PHASE_16 <= _1279;
        else
            if (_72)
                PHASE_16 <= _47;
    end
    assign _1363 = PHASE_16 ? _1362 : _1351;
    assign address_71 = _1548 ? _199 : _1543;
    assign write_enable_71 = _1541 & _1548;
    assign address_72 = _1548 ? _164 : _68;
    assign _1550 = ~ _1548;
    assign read_enable_59 = _1536 & _1550;
    assign _1548 = ~ PHASE_19;
    assign write_enable_72 = _1534 & _1548;
    assign _1552 = write_enable_72 | read_enable_59;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_35
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1552), .regcea(vdd), .wea(write_enable_72), .addra(address_72), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_71), .regceb(vdd), .web(write_enable_71), .addrb(address_71), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1557[131:131]), .sbiterrb(_1557[130:130]), .doutb(_1557[129:66]), .dbiterra(_1557[65:65]), .sbiterra(_1557[64:64]), .douta(_1557[63:0]) );
    assign _1558 = _1557[63:0];
    assign address_73 = PHASE_19 ? _199 : _1543;
    assign _1541 = _129 & _1504;
    assign write_enable_73 = _1541 & PHASE_19;
    assign _1466 = _1458[129:66];
    assign _1465 = _1445[129:66];
    assign _1467 = PHASE_17 ? _1466 : _1465;
    assign _1463 = _1403[129:66];
    assign _1462 = _1389[129:66];
    assign q1_5 = PHASE_18 ? _1463 : _1462;
    assign _1468 = _1370 ? _1467 : q1_5;
    assign address_74 = _1447 ? _1441 : _1440;
    assign _1453 = ~ _1447;
    assign read_enable_60 = _102 & _1453;
    assign address_75 = _1447 ? _60 : _1423;
    assign _1449 = ~ _1447;
    assign read_enable_61 = _102 & _1449;
    assign _1447 = ~ PHASE_17;
    assign write_enable_75 = _1406 & _1447;
    assign _1451 = write_enable_75 | read_enable_61;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_36
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1451), .regcea(vdd), .wea(write_enable_75), .addra(address_75), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_60), .regceb(vdd), .web(write_enable_74), .addrb(address_74), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1458[131:131]), .sbiterrb(_1458[130:130]), .doutb(_1458[129:66]), .dbiterra(_1458[65:65]), .sbiterra(_1458[64:64]), .douta(_1458[63:0]) );
    assign _1459 = _1458[63:0];
    assign _1439 = _172[11:11];
    assign _1438 = _172[10:10];
    assign _1437 = _172[9:9];
    assign _1436 = _172[8:8];
    assign _1435 = _172[7:7];
    assign _1434 = _172[6:6];
    assign _1433 = _172[5:5];
    assign _1432 = _172[4:4];
    assign _1431 = _172[3:3];
    assign _1430 = _172[2:2];
    assign _1429 = _172[1:1];
    assign _1428 = _172[0:0];
    assign _1440 = { _1428, _1429, _1430, _1431, _1432, _1433, _1434, _1435, _1436, _1437, _1438, _1439 };
    assign address_76 = PHASE_17 ? _1441 : _1440;
    assign _1425 = ~ PHASE_17;
    assign read_enable_62 = _102 & _1425;
    assign data_73 = wr_d1;
    assign _1422 = _137[11:11];
    assign _1421 = _137[10:10];
    assign _1420 = _137[9:9];
    assign _1419 = _137[8:8];
    assign _1418 = _137[7:7];
    assign _1417 = _137[6:6];
    assign _1416 = _137[5:5];
    assign _1415 = _137[4:4];
    assign _1414 = _137[3:3];
    assign _1413 = _137[2:2];
    assign _1412 = _137[1:1];
    assign _1411 = _137[0:0];
    assign _1423 = { _1411, _1412, _1413, _1414, _1415, _1416, _1417, _1418, _1419, _1420, _1421, _1422 };
    assign address_77 = PHASE_17 ? _60 : _1423;
    assign _1408 = ~ PHASE_17;
    assign read_enable_63 = _102 & _1408;
    assign _1406 = _62[1:1];
    assign write_enable_77 = _1406 & PHASE_17;
    assign _1410 = write_enable_77 | read_enable_63;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_37
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1410), .regcea(vdd), .wea(write_enable_77), .addra(address_77), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_62), .regceb(vdd), .web(write_enable_76), .addrb(address_76), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1445[131:131]), .sbiterrb(_1445[130:130]), .doutb(_1445[129:66]), .dbiterra(_1445[65:65]), .sbiterra(_1445[64:64]), .douta(_1445[63:0]) );
    assign _1446 = _1445[63:0];
    assign _1367 = ~ PHASE_17;
    assign _51 = _1367;
    always @(posedge _84) begin
        if (_82)
            PHASE_17 <= _1365;
        else
            if (_72)
                PHASE_17 <= _51;
    end
    assign _1460 = PHASE_17 ? _1459 : _1446;
    assign address_78 = _1391 ? _199 : _172;
    assign _1398 = ~ _1391;
    assign read_enable_64 = _102 & _1398;
    assign write_enable_78 = _1382 & _1391;
    assign _1400 = write_enable_78 | read_enable_64;
    assign address_79 = _1391 ? _164 : _137;
    assign _1393 = ~ _1391;
    assign read_enable_65 = _102 & _1393;
    assign _1391 = ~ PHASE_18;
    assign write_enable_79 = _1375 & _1391;
    assign _1395 = write_enable_79 | read_enable_65;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_38
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1395), .regcea(vdd), .wea(write_enable_79), .addra(address_79), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1400), .regceb(vdd), .web(write_enable_78), .addrb(address_78), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1403[131:131]), .sbiterrb(_1403[130:130]), .doutb(_1403[129:66]), .dbiterra(_1403[65:65]), .sbiterra(_1403[64:64]), .douta(_1403[63:0]) );
    assign _1404 = _1403[63:0];
    assign _1471 = _1470[127:64];
    assign data_75 = _1471;
    assign address_80 = PHASE_18 ? _199 : _172;
    assign _1384 = ~ PHASE_18;
    assign read_enable_66 = _102 & _1384;
    assign _1381 = ~ _130;
    assign _1382 = _129 & _1381;
    assign write_enable_80 = _1382 & PHASE_18;
    assign _1386 = write_enable_80 | read_enable_66;
    assign address_81 = PHASE_18 ? _164 : _137;
    assign _1377 = ~ PHASE_18;
    assign read_enable_67 = _102 & _1377;
    assign _1374 = ~ _130;
    assign _1375 = _129 & _1374;
    assign write_enable_81 = _1375 & PHASE_18;
    assign _1379 = write_enable_81 | read_enable_67;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_39
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1379), .regcea(vdd), .wea(write_enable_81), .addra(address_81), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1386), .regceb(vdd), .web(write_enable_80), .addrb(address_80), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1389[131:131]), .sbiterrb(_1389[130:130]), .doutb(_1389[129:66]), .dbiterra(_1389[65:65]), .sbiterra(_1389[64:64]), .douta(_1389[63:0]) );
    assign _1390 = _1389[63:0];
    assign _1472 = ~ PHASE_18;
    assign _53 = _1472;
    always @(posedge _84) begin
        if (_82)
            PHASE_18 <= _1372;
        else
            if (_99)
                PHASE_18 <= _53;
    end
    assign q0_5 = PHASE_18 ? _1404 : _1390;
    always @(posedge _84) begin
        if (_82)
            _1370 <= _1369;
        else
            _1370 <= _92;
    end
    assign _1461 = _1370 ? _1460 : q0_5;
    dp_24
        dp_0
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1461), .d2(_1468), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1470[191:128]), .q2(_1470[127:64]), .q1(_1470[63:0]) );
    assign _1473 = _1470[63:0];
    assign data_79 = _1473;
    assign address_82 = PHASE_19 ? _164 : _68;
    assign _1537 = ~ PHASE_19;
    assign _1536 = _70[1:1];
    assign read_enable_68 = _1536 & _1537;
    always @(posedge _84) begin
        if (_82)
            _1507 <= _1506;
        else
            _1507 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1510 <= _1509;
        else
            _1510 <= _1507;
    end
    always @(posedge _84) begin
        if (_82)
            _1513 <= _1512;
        else
            _1513 <= _1510;
    end
    always @(posedge _84) begin
        if (_82)
            _1516 <= _1515;
        else
            _1516 <= _1513;
    end
    always @(posedge _84) begin
        if (_82)
            _1519 <= _1518;
        else
            _1519 <= _1516;
    end
    always @(posedge _84) begin
        if (_82)
            _1522 <= _1521;
        else
            _1522 <= _1519;
    end
    always @(posedge _84) begin
        if (_82)
            _1525 <= _1524;
        else
            _1525 <= _1522;
    end
    always @(posedge _84) begin
        if (_82)
            _1528 <= _1527;
        else
            _1528 <= _1525;
    end
    always @(posedge _84) begin
        if (_82)
            _1531 <= _1530;
        else
            _1531 <= _1528;
    end
    assign _1532 = ~ _1531;
    always @(posedge _84) begin
        if (_82)
            _1480 <= _1479;
        else
            _1480 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1483 <= _1482;
        else
            _1483 <= _1480;
    end
    always @(posedge _84) begin
        if (_82)
            _1486 <= _1485;
        else
            _1486 <= _1483;
    end
    always @(posedge _84) begin
        if (_82)
            _1489 <= _1488;
        else
            _1489 <= _1486;
    end
    always @(posedge _84) begin
        if (_82)
            _1492 <= _1491;
        else
            _1492 <= _1489;
    end
    always @(posedge _84) begin
        if (_82)
            _1495 <= _1494;
        else
            _1495 <= _1492;
    end
    always @(posedge _84) begin
        if (_82)
            _1498 <= _1497;
        else
            _1498 <= _1495;
    end
    always @(posedge _84) begin
        if (_82)
            _1501 <= _1500;
        else
            _1501 <= _1498;
    end
    always @(posedge _84) begin
        if (_82)
            _1504 <= _1503;
        else
            _1504 <= _1501;
    end
    assign _1533 = _1504 & _1532;
    assign _1534 = _129 & _1533;
    assign write_enable_82 = _1534 & PHASE_19;
    assign _1539 = write_enable_82 | read_enable_68;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_40
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1539), .regcea(vdd), .wea(write_enable_82), .addra(address_82), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_73), .regceb(vdd), .web(write_enable_73), .addrb(address_73), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1546[131:131]), .sbiterrb(_1546[130:130]), .doutb(_1546[129:66]), .dbiterra(_1546[65:65]), .sbiterra(_1546[64:64]), .douta(_1546[63:0]) );
    assign _1547 = _1546[63:0];
    assign _1477 = ~ PHASE_19;
    assign _55 = _1477;
    always @(posedge _84) begin
        if (_82)
            PHASE_19 <= _1475;
        else
            if (_72)
                PHASE_19 <= _55;
    end
    assign _1559 = PHASE_19 ? _1558 : _1547;
    assign address_83 = _1744 ? _199 : _1739;
    assign write_enable_83 = _1737 & _1744;
    assign address_84 = _1744 ? _164 : _68;
    assign _1746 = ~ _1744;
    assign read_enable_69 = _1732 & _1746;
    assign _1744 = ~ PHASE_22;
    assign write_enable_84 = _1730 & _1744;
    assign _1748 = write_enable_84 | read_enable_69;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_41
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1748), .regcea(vdd), .wea(write_enable_84), .addra(address_84), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_83), .regceb(vdd), .web(write_enable_83), .addrb(address_83), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1753[131:131]), .sbiterrb(_1753[130:130]), .doutb(_1753[129:66]), .dbiterra(_1753[65:65]), .sbiterra(_1753[64:64]), .douta(_1753[63:0]) );
    assign _1754 = _1753[63:0];
    assign address_85 = PHASE_22 ? _199 : _1739;
    assign _1737 = _129 & _1700;
    assign write_enable_85 = _1737 & PHASE_22;
    assign _292 = _91[521:518];
    assign _291 = _91[517:517];
    assign _289 = _91[513:513];
    assign _288 = _91[512:449];
    assign _287 = _91[448:385];
    assign _286 = _91[384:321];
    assign _285 = _91[320:257];
    assign _284 = _91[256:193];
    assign _283 = _91[192:129];
    assign _282 = _91[128:65];
    assign _1662 = _1654[129:66];
    assign _1661 = _1641[129:66];
    assign _1663 = PHASE_20 ? _1662 : _1661;
    assign _1659 = _1599[129:66];
    assign _1658 = _1585[129:66];
    assign q1_6 = PHASE_21 ? _1659 : _1658;
    assign _1664 = _1566 ? _1663 : q1_6;
    assign address_86 = _1643 ? _1637 : _1636;
    assign _1649 = ~ _1643;
    assign read_enable_70 = _102 & _1649;
    assign address_87 = _1643 ? _60 : _1619;
    assign _1645 = ~ _1643;
    assign read_enable_71 = _102 & _1645;
    assign _1643 = ~ PHASE_20;
    assign write_enable_87 = _1602 & _1643;
    assign _1647 = write_enable_87 | read_enable_71;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_42
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1647), .regcea(vdd), .wea(write_enable_87), .addra(address_87), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_70), .regceb(vdd), .web(write_enable_86), .addrb(address_86), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1654[131:131]), .sbiterrb(_1654[130:130]), .doutb(_1654[129:66]), .dbiterra(_1654[65:65]), .sbiterra(_1654[64:64]), .douta(_1654[63:0]) );
    assign _1655 = _1654[63:0];
    assign _1635 = _172[11:11];
    assign _1634 = _172[10:10];
    assign _1633 = _172[9:9];
    assign _1632 = _172[8:8];
    assign _1631 = _172[7:7];
    assign _1630 = _172[6:6];
    assign _1629 = _172[5:5];
    assign _1628 = _172[4:4];
    assign _1627 = _172[3:3];
    assign _1626 = _172[2:2];
    assign _1625 = _172[1:1];
    assign _1624 = _172[0:0];
    assign _1636 = { _1624, _1625, _1626, _1627, _1628, _1629, _1630, _1631, _1632, _1633, _1634, _1635 };
    assign address_88 = PHASE_20 ? _1637 : _1636;
    assign _1621 = ~ PHASE_20;
    assign read_enable_72 = _102 & _1621;
    assign data_85 = wr_d0;
    assign _60 = wr_addr;
    assign _1618 = _137[11:11];
    assign _1617 = _137[10:10];
    assign _1616 = _137[9:9];
    assign _1615 = _137[8:8];
    assign _1614 = _137[7:7];
    assign _1613 = _137[6:6];
    assign _1612 = _137[5:5];
    assign _1611 = _137[4:4];
    assign _1610 = _137[3:3];
    assign _1609 = _137[2:2];
    assign _1608 = _137[1:1];
    assign _1607 = _137[0:0];
    assign _1619 = { _1607, _1608, _1609, _1610, _1611, _1612, _1613, _1614, _1615, _1616, _1617, _1618 };
    assign address_89 = PHASE_20 ? _60 : _1619;
    assign _1604 = ~ PHASE_20;
    assign read_enable_73 = _102 & _1604;
    assign _62 = wr_en;
    assign _1602 = _62[0:0];
    assign write_enable_89 = _1602 & PHASE_20;
    assign _1606 = write_enable_89 | read_enable_73;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_43
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1606), .regcea(vdd), .wea(write_enable_89), .addra(address_89), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_72), .regceb(vdd), .web(write_enable_88), .addrb(address_88), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1641[131:131]), .sbiterrb(_1641[130:130]), .doutb(_1641[129:66]), .dbiterra(_1641[65:65]), .sbiterra(_1641[64:64]), .douta(_1641[63:0]) );
    assign _1642 = _1641[63:0];
    assign _1563 = ~ PHASE_20;
    assign _63 = _1563;
    always @(posedge _84) begin
        if (_82)
            PHASE_20 <= _1561;
        else
            if (_72)
                PHASE_20 <= _63;
    end
    assign _1656 = PHASE_20 ? _1655 : _1642;
    assign address_90 = _1587 ? _199 : _172;
    assign _1594 = ~ _1587;
    assign read_enable_74 = _102 & _1594;
    assign write_enable_90 = _1578 & _1587;
    assign _1596 = write_enable_90 | read_enable_74;
    assign address_91 = _1587 ? _164 : _137;
    assign _1589 = ~ _1587;
    assign read_enable_75 = _102 & _1589;
    assign _1587 = ~ PHASE_21;
    assign write_enable_91 = _1571 & _1587;
    assign _1591 = write_enable_91 | read_enable_75;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_44
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1591), .regcea(vdd), .wea(write_enable_91), .addra(address_91), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1596), .regceb(vdd), .web(write_enable_90), .addrb(address_90), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1599[131:131]), .sbiterrb(_1599[130:130]), .doutb(_1599[129:66]), .dbiterra(_1599[65:65]), .sbiterra(_1599[64:64]), .douta(_1599[63:0]) );
    assign _1600 = _1599[63:0];
    assign _1667 = _1666[127:64];
    assign data_87 = _1667;
    always @(posedge _84) begin
        if (_82)
            _175 <= _174;
        else
            _175 <= _172;
    end
    always @(posedge _84) begin
        if (_82)
            _178 <= _177;
        else
            _178 <= _175;
    end
    always @(posedge _84) begin
        if (_82)
            _181 <= _180;
        else
            _181 <= _178;
    end
    always @(posedge _84) begin
        if (_82)
            _184 <= _183;
        else
            _184 <= _181;
    end
    always @(posedge _84) begin
        if (_82)
            _187 <= _186;
        else
            _187 <= _184;
    end
    always @(posedge _84) begin
        if (_82)
            _190 <= _189;
        else
            _190 <= _187;
    end
    always @(posedge _84) begin
        if (_82)
            _193 <= _192;
        else
            _193 <= _190;
    end
    always @(posedge _84) begin
        if (_82)
            _196 <= _195;
        else
            _196 <= _193;
    end
    always @(posedge _84) begin
        if (_82)
            _199 <= _198;
        else
            _199 <= _196;
    end
    assign _172 = _91[64:53];
    assign address_92 = PHASE_21 ? _199 : _172;
    assign _1580 = ~ PHASE_21;
    assign read_enable_76 = _102 & _1580;
    assign _1577 = ~ _130;
    assign _1578 = _129 & _1577;
    assign write_enable_92 = _1578 & PHASE_21;
    assign _1582 = write_enable_92 | read_enable_76;
    assign address_93 = PHASE_21 ? _164 : _137;
    assign _1573 = ~ PHASE_21;
    assign read_enable_77 = _102 & _1573;
    assign _1570 = ~ _130;
    assign _1571 = _129 & _1570;
    assign write_enable_93 = _1571 & PHASE_21;
    assign _1575 = write_enable_93 | read_enable_77;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_45
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1575), .regcea(vdd), .wea(write_enable_93), .addra(address_93), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1582), .regceb(vdd), .web(write_enable_92), .addrb(address_92), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1585[131:131]), .sbiterrb(_1585[130:130]), .doutb(_1585[129:66]), .dbiterra(_1585[65:65]), .sbiterra(_1585[64:64]), .douta(_1585[63:0]) );
    assign _1586 = _1585[63:0];
    assign _99 = _91[523:523];
    assign _1668 = ~ PHASE_21;
    assign _65 = _1668;
    always @(posedge _84) begin
        if (_82)
            PHASE_21 <= _1568;
        else
            if (_99)
                PHASE_21 <= _65;
    end
    assign q0_6 = PHASE_21 ? _1600 : _1586;
    assign _92 = _91[514:514];
    always @(posedge _84) begin
        if (_82)
            _1566 <= _1565;
        else
            _1566 <= _92;
    end
    assign _1657 = _1566 ? _1656 : q0_6;
    dp_23
        dp
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1657), .d2(_1664), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1666[191:128]), .q2(_1666[127:64]), .q1(_1666[63:0]) );
    assign _1669 = _1666[63:0];
    assign data_91 = _1669;
    assign _137 = _91[52:41];
    always @(posedge _84) begin
        if (_82)
            _140 <= _139;
        else
            _140 <= _137;
    end
    always @(posedge _84) begin
        if (_82)
            _143 <= _142;
        else
            _143 <= _140;
    end
    always @(posedge _84) begin
        if (_82)
            _146 <= _145;
        else
            _146 <= _143;
    end
    always @(posedge _84) begin
        if (_82)
            _149 <= _148;
        else
            _149 <= _146;
    end
    always @(posedge _84) begin
        if (_82)
            _152 <= _151;
        else
            _152 <= _149;
    end
    always @(posedge _84) begin
        if (_82)
            _155 <= _154;
        else
            _155 <= _152;
    end
    always @(posedge _84) begin
        if (_82)
            _158 <= _157;
        else
            _158 <= _155;
    end
    always @(posedge _84) begin
        if (_82)
            _161 <= _160;
        else
            _161 <= _158;
    end
    always @(posedge _84) begin
        if (_82)
            _164 <= _163;
        else
            _164 <= _161;
    end
    assign _68 = rd_addr;
    assign address_94 = PHASE_22 ? _164 : _68;
    assign _1733 = ~ PHASE_22;
    assign _70 = rd_en;
    assign _1732 = _70[0:0];
    assign read_enable_78 = _1732 & _1733;
    assign _290 = _91[516:516];
    always @(posedge _84) begin
        if (_82)
            _1703 <= _1702;
        else
            _1703 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1706 <= _1705;
        else
            _1706 <= _1703;
    end
    always @(posedge _84) begin
        if (_82)
            _1709 <= _1708;
        else
            _1709 <= _1706;
    end
    always @(posedge _84) begin
        if (_82)
            _1712 <= _1711;
        else
            _1712 <= _1709;
    end
    always @(posedge _84) begin
        if (_82)
            _1715 <= _1714;
        else
            _1715 <= _1712;
    end
    always @(posedge _84) begin
        if (_82)
            _1718 <= _1717;
        else
            _1718 <= _1715;
    end
    always @(posedge _84) begin
        if (_82)
            _1721 <= _1720;
        else
            _1721 <= _1718;
    end
    always @(posedge _84) begin
        if (_82)
            _1724 <= _1723;
        else
            _1724 <= _1721;
    end
    always @(posedge _84) begin
        if (_82)
            _1727 <= _1726;
        else
            _1727 <= _1724;
    end
    assign _1728 = ~ _1727;
    assign _130 = _91[515:515];
    always @(posedge _84) begin
        if (_82)
            _1676 <= _1675;
        else
            _1676 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1679 <= _1678;
        else
            _1679 <= _1676;
    end
    always @(posedge _84) begin
        if (_82)
            _1682 <= _1681;
        else
            _1682 <= _1679;
    end
    always @(posedge _84) begin
        if (_82)
            _1685 <= _1684;
        else
            _1685 <= _1682;
    end
    always @(posedge _84) begin
        if (_82)
            _1688 <= _1687;
        else
            _1688 <= _1685;
    end
    always @(posedge _84) begin
        if (_82)
            _1691 <= _1690;
        else
            _1691 <= _1688;
    end
    always @(posedge _84) begin
        if (_82)
            _1694 <= _1693;
        else
            _1694 <= _1691;
    end
    always @(posedge _84) begin
        if (_82)
            _1697 <= _1696;
        else
            _1697 <= _1694;
    end
    always @(posedge _84) begin
        if (_82)
            _1700 <= _1699;
        else
            _1700 <= _1697;
    end
    assign _1729 = _1700 & _1728;
    assign _102 = _91[522:522];
    always @(posedge _84) begin
        if (_82)
            _105 <= _104;
        else
            _105 <= _102;
    end
    always @(posedge _84) begin
        if (_82)
            _108 <= _107;
        else
            _108 <= _105;
    end
    always @(posedge _84) begin
        if (_82)
            _111 <= _110;
        else
            _111 <= _108;
    end
    always @(posedge _84) begin
        if (_82)
            _114 <= _113;
        else
            _114 <= _111;
    end
    always @(posedge _84) begin
        if (_82)
            _117 <= _116;
        else
            _117 <= _114;
    end
    always @(posedge _84) begin
        if (_82)
            _120 <= _119;
        else
            _120 <= _117;
    end
    always @(posedge _84) begin
        if (_82)
            _123 <= _122;
        else
            _123 <= _120;
    end
    always @(posedge _84) begin
        if (_82)
            _126 <= _125;
        else
            _126 <= _123;
    end
    always @(posedge _84) begin
        if (_82)
            _129 <= _128;
        else
            _129 <= _126;
    end
    assign _1730 = _129 & _1729;
    assign write_enable_94 = _1730 & PHASE_22;
    assign _1735 = write_enable_94 | read_enable_78;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_46
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1735), .regcea(vdd), .wea(write_enable_94), .addra(address_94), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_85), .regceb(vdd), .web(write_enable_85), .addrb(address_85), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1742[131:131]), .sbiterrb(_1742[130:130]), .doutb(_1742[129:66]), .dbiterra(_1742[65:65]), .sbiterra(_1742[64:64]), .douta(_1742[63:0]) );
    assign _1743 = _1742[63:0];
    assign _72 = flip;
    assign _1673 = ~ PHASE_22;
    assign _73 = _1673;
    always @(posedge _84) begin
        if (_82)
            PHASE_22 <= _1671;
        else
            if (_72)
                PHASE_22 <= _73;
    end
    assign _1755 = PHASE_22 ? _1754 : _1743;
    assign _76 = first_4step_pass;
    assign _78 = first_iter;
    assign _80 = start;
    assign _82 = clear;
    assign _84 = clock;
    ctrl
        ctrl
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .first_4step_pass(_76), .flip(_91[523:523]), .read_write_enable(_91[522:522]), .index(_91[521:518]), .valid(_91[517:517]), .twiddle_stage(_91[516:516]), .last_stage(_91[515:515]), .first_stage(_91[514:514]), .start_twiddles(_91[513:513]), .omegas6(_91[512:449]), .omegas5(_91[448:385]), .omegas4(_91[384:321]), .omegas3(_91[320:257]), .omegas2(_91[256:193]), .omegas1(_91[192:129]), .omegas0(_91[128:65]), .addr2(_91[64:53]), .addr1(_91[52:41]), .m(_91[40:29]), .k(_91[28:17]), .j(_91[16:5]), .i(_91[4:1]), .done_(_91[0:0]) );
    assign _1756 = _91[0:0];

    /* aliases */
    assign data_0 = data;
    assign data_2 = data_1;
    assign data_4 = data_3;
    assign data_5 = data_3;
    assign data_6 = data_3;
    assign data_8 = data_7;
    assign data_9 = data_7;
    assign data_10 = data_7;
    assign data_12 = data_11;
    assign data_14 = data_13;
    assign data_16 = data_15;
    assign data_17 = data_15;
    assign data_18 = data_15;
    assign data_20 = data_19;
    assign data_21 = data_19;
    assign data_22 = data_19;
    assign data_24 = data_23;
    assign data_26 = data_25;
    assign data_28 = data_27;
    assign data_29 = data_27;
    assign data_30 = data_27;
    assign data_32 = data_31;
    assign data_33 = data_31;
    assign data_34 = data_31;
    assign data_36 = data_35;
    assign data_38 = data_37;
    assign data_40 = data_39;
    assign data_41 = data_39;
    assign data_42 = data_39;
    assign data_44 = data_43;
    assign data_45 = data_43;
    assign data_46 = data_43;
    assign data_48 = data_47;
    assign data_50 = data_49;
    assign data_52 = data_51;
    assign data_53 = data_51;
    assign data_54 = data_51;
    assign data_56 = data_55;
    assign data_57 = data_55;
    assign data_58 = data_55;
    assign data_60 = data_59;
    assign data_62 = data_61;
    assign data_64 = data_63;
    assign data_65 = data_63;
    assign data_66 = data_63;
    assign data_68 = data_67;
    assign data_69 = data_67;
    assign data_70 = data_67;
    assign data_72 = data_71;
    assign data_74 = data_73;
    assign data_76 = data_75;
    assign data_77 = data_75;
    assign data_78 = data_75;
    assign data_80 = data_79;
    assign data_81 = data_79;
    assign data_82 = data_79;
    assign data_84 = data_83;
    assign data_86 = data_85;
    assign data_88 = data_87;
    assign data_89 = data_87;
    assign data_90 = data_87;
    assign data_92 = data_91;
    assign data_93 = data_91;
    assign data_94 = data_91;

    /* output assignments */
    assign done_ = _1756;
    assign rd_q0 = _1755;
    assign rd_q1 = _1559;
    assign rd_q2 = _1363;
    assign rd_q3 = _1167;
    assign rd_q4 = _971;
    assign rd_q5 = _775;
    assign rd_q6 = _579;
    assign rd_q7 = _383;

endmodule
module dp_31 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0111100010011001111011110010110000010101011010110010100000110001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0100010101011101011101010011001111101010110011010001000101010111;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0110100110010111111010001101100011001001101111010100100000100101;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1111101111010100000111000110101110001100101010100011001100000010;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_32 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0001100001101001111110100111111110111000110010000010011011110100;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1111110001000101101010101010100100111100101011011000000100111100;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0100001010110000001101000000101010000000011110111001101000111101;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0100011111101001000011110000001000111010101011110101010100100101;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1100111011101001001111010011000100010100101000011000000011000111;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0110100101101111110010001001101110011101101001011110000011100001;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1100001001011111000111001110000000001100100011011001101101100111;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_33 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1000010000100010101000000000111110001110011111011110010000111111;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0000101111001000100000001011001110110011001101111111011010000101;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0011110010111001010110011011000110010111010110100011001100100111;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1111100101010101101110010000101110110010011010100110000011000000;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0111111010110111000101110011011011100010101100111010000100000110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1001110001100101101001000011100011101100100110101001011111111000;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0110101111000000010111100100011101010101010001100110100011000010;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_34 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1101011010101010101100111101101011101110011110100000110011000011;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0011110101010010010000101110111110001011011110110110010010111001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1000001101101101010001010010111001000010111000101011100011100110;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1000000000010101010101101101000101010110000010111110001110111000;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0101110100110000000100110101011101000010111111000111010000001011;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1100001011100100110011000100001001100010000010000101000110100011;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0111110011001000110011000001001011011101111010111000111010000010;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_35 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0011000101111100111000111101000110001100011110101101101000010101;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1010001101101010010111100101011111010001100010010100010001010001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1010101100000000110010110011010110110001111111010100000010011110;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0011110101010110000000001101011100010100100101111100001010111100;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0001001000111000010111110001101011011001000001111111010110000000;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0000000110011111011011110111001101111001110110010011010011110001;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0110110010110000111011001100000000010111101011101101100010111100;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_36 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0000011101101001011001000000101010000101001000001111110101011110;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1100110000010111010111000011011111001001110111110101100110110100;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0011110000011000000100100001110101111011111111000001000100111010;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1000101010110100010111011000000010111011100001101001011001101111;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1110001110011100011000011110000101011111101011100011110010100110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1110111100010111011111001000000001011100101111111101111110000101;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0101100010111110011100110111001111001001000001011110110110110010;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_37 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0101000111001001010010110111011001100011110011111111110010111001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0111001111011001100001101101101110110111101001010001010011001101;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1010000001111100110100111101111011010101010101110110100000101110;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0110100110111100001101111100000111000010011011001010010111000011;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1100100010110010000000011011001100000010111000101000000110010110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0100100010101101111000110100110001111001100110001001111000111111;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1011001111101011010100101110010011000101101010010001011100000111;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_38 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1100000001010000000100100000100111101111010000100000001100000011;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0001110000000100101011001111001110000101010001000100111011101111;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0110000101101100010100011110001010010011011010101000000000100111;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0110101010010110110001001110100010101101100101010001110111001100;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0101000010000011110011000110111011011100001001000011111000110001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0010111110010100110000110000001100100101110011011100011011100111;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0001001110110001100110001111101111010100011111111100000011111001;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module parallel_cores_3 (
    wr_d7,
    wr_d6,
    wr_d5,
    wr_d4,
    wr_d3,
    wr_d2,
    wr_d1,
    wr_d0,
    wr_addr,
    wr_en,
    rd_addr,
    rd_en,
    flip,
    first_4step_pass,
    first_iter,
    start,
    clear,
    clock,
    done_,
    rd_q0,
    rd_q1,
    rd_q2,
    rd_q3,
    rd_q4,
    rd_q5,
    rd_q6,
    rd_q7
);

    input [63:0] wr_d7;
    input [63:0] wr_d6;
    input [63:0] wr_d5;
    input [63:0] wr_d4;
    input [63:0] wr_d3;
    input [63:0] wr_d2;
    input [63:0] wr_d1;
    input [63:0] wr_d0;
    input [11:0] wr_addr;
    input [7:0] wr_en;
    input [11:0] rd_addr;
    input [7:0] rd_en;
    input flip;
    input first_4step_pass;
    input first_iter;
    input start;
    input clear;
    input clock;
    output done_;
    output [63:0] rd_q0;
    output [63:0] rd_q1;
    output [63:0] rd_q2;
    output [63:0] rd_q3;
    output [63:0] rd_q4;
    output [63:0] rd_q5;
    output [63:0] rd_q6;
    output [63:0] rd_q7;

    /* signal declarations */
    wire [11:0] address;
    wire write_enable;
    wire [11:0] address_0;
    wire _374;
    wire read_enable;
    wire _372;
    wire write_enable_0;
    wire _376;
    wire [131:0] _381;
    wire [63:0] _382;
    wire [11:0] _367 = 12'b000000000000;
    wire [11:0] address_1;
    wire _365;
    wire write_enable_1;
    wire [63:0] _279;
    wire [63:0] _278;
    wire [63:0] _280;
    wire [63:0] _276;
    wire [63:0] _275;
    wire [63:0] q1;
    wire [63:0] _281;
    wire [11:0] address_2;
    wire write_enable_2 = 1'b0;
    wire _266;
    wire read_enable_0;
    wire [11:0] address_3;
    wire _262;
    wire read_enable_1;
    wire _260;
    wire write_enable_3;
    wire _264;
    wire [131:0] _271;
    wire [63:0] _272;
    wire [63:0] data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_0;
    wire [11:0] _254 = 12'b000000000000;
    wire _252;
    wire _251;
    wire _250;
    wire _249;
    wire _248;
    wire _247;
    wire _246;
    wire _245;
    wire _244;
    wire _243;
    wire _242;
    wire _241;
    wire [11:0] _253;
    wire [11:0] address_4;
    wire write_enable_4 = 1'b0;
    wire _238;
    wire read_enable_2;
    wire [63:0] data_1;
    wire [63:0] data_2;
    wire _235;
    wire _234;
    wire _233;
    wire _232;
    wire _231;
    wire _230;
    wire _229;
    wire _228;
    wire _227;
    wire _226;
    wire _225;
    wire _224;
    wire [11:0] _236;
    wire [11:0] address_5;
    wire _221;
    wire read_enable_3;
    wire _219;
    wire write_enable_5;
    wire _223;
    wire [131:0] _258;
    wire [63:0] _259;
    wire _87 = 1'b0;
    wire _86 = 1'b0;
    wire _89;
    wire _3;
    reg PHASE;
    wire [63:0] _273;
    wire [11:0] address_6;
    wire _211;
    wire read_enable_4;
    wire write_enable_6;
    wire _213;
    wire [11:0] address_7;
    wire _206;
    wire read_enable_5;
    wire _204;
    wire write_enable_7;
    wire _208;
    wire [131:0] _216;
    wire [63:0] _217;
    wire [63:0] _295;
    wire [63:0] data_3;
    wire [63:0] data_4;
    wire [63:0] data_5;
    wire [63:0] data_6;
    wire [11:0] address_8;
    wire _169;
    wire read_enable_6;
    wire _166;
    wire _167;
    wire write_enable_8;
    wire _171;
    wire [11:0] address_9;
    wire _134;
    wire read_enable_7;
    wire _131;
    wire _132;
    wire write_enable_9;
    wire _136;
    wire [131:0] _202;
    wire [63:0] _203;
    wire _98 = 1'b0;
    wire _97 = 1'b0;
    wire _296;
    wire _5;
    reg PHASE_0;
    wire [63:0] q0;
    wire _94 = 1'b0;
    wire _93 = 1'b0;
    reg _96;
    wire [63:0] _274;
    wire [191:0] _294;
    wire [63:0] _297;
    wire [63:0] data_7;
    wire [63:0] data_8;
    wire [63:0] data_9;
    wire [63:0] data_10;
    wire [11:0] address_10;
    wire _361;
    wire _360;
    wire read_enable_8;
    wire _354 = 1'b0;
    wire _353 = 1'b0;
    wire _351 = 1'b0;
    wire _350 = 1'b0;
    wire _348 = 1'b0;
    wire _347 = 1'b0;
    wire _345 = 1'b0;
    wire _344 = 1'b0;
    wire _342 = 1'b0;
    wire _341 = 1'b0;
    wire _339 = 1'b0;
    wire _338 = 1'b0;
    wire _336 = 1'b0;
    wire _335 = 1'b0;
    wire _333 = 1'b0;
    wire _332 = 1'b0;
    wire _330 = 1'b0;
    wire _329 = 1'b0;
    reg _331;
    reg _334;
    reg _337;
    reg _340;
    reg _343;
    reg _346;
    reg _349;
    reg _352;
    reg _355;
    wire _356;
    wire _327 = 1'b0;
    wire _326 = 1'b0;
    wire _324 = 1'b0;
    wire _323 = 1'b0;
    wire _321 = 1'b0;
    wire _320 = 1'b0;
    wire _318 = 1'b0;
    wire _317 = 1'b0;
    wire _315 = 1'b0;
    wire _314 = 1'b0;
    wire _312 = 1'b0;
    wire _311 = 1'b0;
    wire _309 = 1'b0;
    wire _308 = 1'b0;
    wire _306 = 1'b0;
    wire _305 = 1'b0;
    wire _303 = 1'b0;
    wire _302 = 1'b0;
    reg _304;
    reg _307;
    reg _310;
    reg _313;
    reg _316;
    reg _319;
    reg _322;
    reg _325;
    reg _328;
    wire _357;
    wire _358;
    wire write_enable_10;
    wire _363;
    wire [131:0] _370;
    wire [63:0] _371;
    wire _299 = 1'b0;
    wire _298 = 1'b0;
    wire _301;
    wire _7;
    reg PHASE_1;
    wire [63:0] _383;
    wire [11:0] address_11;
    wire write_enable_11;
    wire [11:0] address_12;
    wire _570;
    wire read_enable_9;
    wire _568;
    wire write_enable_12;
    wire _572;
    wire [131:0] _577;
    wire [63:0] _578;
    wire [11:0] _563 = 12'b000000000000;
    wire [11:0] address_13;
    wire _561;
    wire write_enable_13;
    wire [63:0] _486;
    wire [63:0] _485;
    wire [63:0] _487;
    wire [63:0] _483;
    wire [63:0] _482;
    wire [63:0] q1_0;
    wire [63:0] _488;
    wire [11:0] address_14;
    wire write_enable_14 = 1'b0;
    wire _473;
    wire read_enable_10;
    wire [11:0] address_15;
    wire _469;
    wire read_enable_11;
    wire _467;
    wire write_enable_15;
    wire _471;
    wire [131:0] _478;
    wire [63:0] _479;
    wire [63:0] data_11 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_12;
    wire [11:0] _461 = 12'b000000000000;
    wire _459;
    wire _458;
    wire _457;
    wire _456;
    wire _455;
    wire _454;
    wire _453;
    wire _452;
    wire _451;
    wire _450;
    wire _449;
    wire _448;
    wire [11:0] _460;
    wire [11:0] address_16;
    wire write_enable_16 = 1'b0;
    wire _445;
    wire read_enable_12;
    wire [63:0] data_13;
    wire [63:0] data_14;
    wire _442;
    wire _441;
    wire _440;
    wire _439;
    wire _438;
    wire _437;
    wire _436;
    wire _435;
    wire _434;
    wire _433;
    wire _432;
    wire _431;
    wire [11:0] _443;
    wire [11:0] address_17;
    wire _428;
    wire read_enable_13;
    wire _426;
    wire write_enable_17;
    wire _430;
    wire [131:0] _465;
    wire [63:0] _466;
    wire _385 = 1'b0;
    wire _384 = 1'b0;
    wire _387;
    wire _11;
    reg PHASE_2;
    wire [63:0] _480;
    wire [11:0] address_18;
    wire _418;
    wire read_enable_14;
    wire write_enable_18;
    wire _420;
    wire [11:0] address_19;
    wire _413;
    wire read_enable_15;
    wire _411;
    wire write_enable_19;
    wire _415;
    wire [131:0] _423;
    wire [63:0] _424;
    wire [63:0] _491;
    wire [63:0] data_15;
    wire [63:0] data_16;
    wire [63:0] data_17;
    wire [63:0] data_18;
    wire [11:0] address_20;
    wire _404;
    wire read_enable_16;
    wire _401;
    wire _402;
    wire write_enable_20;
    wire _406;
    wire [11:0] address_21;
    wire _397;
    wire read_enable_17;
    wire _394;
    wire _395;
    wire write_enable_21;
    wire _399;
    wire [131:0] _409;
    wire [63:0] _410;
    wire _392 = 1'b0;
    wire _391 = 1'b0;
    wire _492;
    wire _13;
    reg PHASE_3;
    wire [63:0] q0_0;
    wire _389 = 1'b0;
    wire _388 = 1'b0;
    reg _390;
    wire [63:0] _481;
    wire [191:0] _490;
    wire [63:0] _493;
    wire [63:0] data_19;
    wire [63:0] data_20;
    wire [63:0] data_21;
    wire [63:0] data_22;
    wire [11:0] address_22;
    wire _557;
    wire _556;
    wire read_enable_18;
    wire _550 = 1'b0;
    wire _549 = 1'b0;
    wire _547 = 1'b0;
    wire _546 = 1'b0;
    wire _544 = 1'b0;
    wire _543 = 1'b0;
    wire _541 = 1'b0;
    wire _540 = 1'b0;
    wire _538 = 1'b0;
    wire _537 = 1'b0;
    wire _535 = 1'b0;
    wire _534 = 1'b0;
    wire _532 = 1'b0;
    wire _531 = 1'b0;
    wire _529 = 1'b0;
    wire _528 = 1'b0;
    wire _526 = 1'b0;
    wire _525 = 1'b0;
    reg _527;
    reg _530;
    reg _533;
    reg _536;
    reg _539;
    reg _542;
    reg _545;
    reg _548;
    reg _551;
    wire _552;
    wire _523 = 1'b0;
    wire _522 = 1'b0;
    wire _520 = 1'b0;
    wire _519 = 1'b0;
    wire _517 = 1'b0;
    wire _516 = 1'b0;
    wire _514 = 1'b0;
    wire _513 = 1'b0;
    wire _511 = 1'b0;
    wire _510 = 1'b0;
    wire _508 = 1'b0;
    wire _507 = 1'b0;
    wire _505 = 1'b0;
    wire _504 = 1'b0;
    wire _502 = 1'b0;
    wire _501 = 1'b0;
    wire _499 = 1'b0;
    wire _498 = 1'b0;
    reg _500;
    reg _503;
    reg _506;
    reg _509;
    reg _512;
    reg _515;
    reg _518;
    reg _521;
    reg _524;
    wire _553;
    wire _554;
    wire write_enable_22;
    wire _559;
    wire [131:0] _566;
    wire [63:0] _567;
    wire _495 = 1'b0;
    wire _494 = 1'b0;
    wire _497;
    wire _15;
    reg PHASE_4;
    wire [63:0] _579;
    wire [11:0] address_23;
    wire write_enable_23;
    wire [11:0] address_24;
    wire _766;
    wire read_enable_19;
    wire _764;
    wire write_enable_24;
    wire _768;
    wire [131:0] _773;
    wire [63:0] _774;
    wire [11:0] _759 = 12'b000000000000;
    wire [11:0] address_25;
    wire _757;
    wire write_enable_25;
    wire [63:0] _682;
    wire [63:0] _681;
    wire [63:0] _683;
    wire [63:0] _679;
    wire [63:0] _678;
    wire [63:0] q1_1;
    wire [63:0] _684;
    wire [11:0] address_26;
    wire write_enable_26 = 1'b0;
    wire _669;
    wire read_enable_20;
    wire [11:0] address_27;
    wire _665;
    wire read_enable_21;
    wire _663;
    wire write_enable_27;
    wire _667;
    wire [131:0] _674;
    wire [63:0] _675;
    wire [63:0] data_23 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_24;
    wire [11:0] _657 = 12'b000000000000;
    wire _655;
    wire _654;
    wire _653;
    wire _652;
    wire _651;
    wire _650;
    wire _649;
    wire _648;
    wire _647;
    wire _646;
    wire _645;
    wire _644;
    wire [11:0] _656;
    wire [11:0] address_28;
    wire write_enable_28 = 1'b0;
    wire _641;
    wire read_enable_22;
    wire [63:0] data_25;
    wire [63:0] data_26;
    wire _638;
    wire _637;
    wire _636;
    wire _635;
    wire _634;
    wire _633;
    wire _632;
    wire _631;
    wire _630;
    wire _629;
    wire _628;
    wire _627;
    wire [11:0] _639;
    wire [11:0] address_29;
    wire _624;
    wire read_enable_23;
    wire _622;
    wire write_enable_29;
    wire _626;
    wire [131:0] _661;
    wire [63:0] _662;
    wire _581 = 1'b0;
    wire _580 = 1'b0;
    wire _583;
    wire _19;
    reg PHASE_5;
    wire [63:0] _676;
    wire [11:0] address_30;
    wire _614;
    wire read_enable_24;
    wire write_enable_30;
    wire _616;
    wire [11:0] address_31;
    wire _609;
    wire read_enable_25;
    wire _607;
    wire write_enable_31;
    wire _611;
    wire [131:0] _619;
    wire [63:0] _620;
    wire [63:0] _687;
    wire [63:0] data_27;
    wire [63:0] data_28;
    wire [63:0] data_29;
    wire [63:0] data_30;
    wire [11:0] address_32;
    wire _600;
    wire read_enable_26;
    wire _597;
    wire _598;
    wire write_enable_32;
    wire _602;
    wire [11:0] address_33;
    wire _593;
    wire read_enable_27;
    wire _590;
    wire _591;
    wire write_enable_33;
    wire _595;
    wire [131:0] _605;
    wire [63:0] _606;
    wire _588 = 1'b0;
    wire _587 = 1'b0;
    wire _688;
    wire _21;
    reg PHASE_6;
    wire [63:0] q0_1;
    wire _585 = 1'b0;
    wire _584 = 1'b0;
    reg _586;
    wire [63:0] _677;
    wire [191:0] _686;
    wire [63:0] _689;
    wire [63:0] data_31;
    wire [63:0] data_32;
    wire [63:0] data_33;
    wire [63:0] data_34;
    wire [11:0] address_34;
    wire _753;
    wire _752;
    wire read_enable_28;
    wire _746 = 1'b0;
    wire _745 = 1'b0;
    wire _743 = 1'b0;
    wire _742 = 1'b0;
    wire _740 = 1'b0;
    wire _739 = 1'b0;
    wire _737 = 1'b0;
    wire _736 = 1'b0;
    wire _734 = 1'b0;
    wire _733 = 1'b0;
    wire _731 = 1'b0;
    wire _730 = 1'b0;
    wire _728 = 1'b0;
    wire _727 = 1'b0;
    wire _725 = 1'b0;
    wire _724 = 1'b0;
    wire _722 = 1'b0;
    wire _721 = 1'b0;
    reg _723;
    reg _726;
    reg _729;
    reg _732;
    reg _735;
    reg _738;
    reg _741;
    reg _744;
    reg _747;
    wire _748;
    wire _719 = 1'b0;
    wire _718 = 1'b0;
    wire _716 = 1'b0;
    wire _715 = 1'b0;
    wire _713 = 1'b0;
    wire _712 = 1'b0;
    wire _710 = 1'b0;
    wire _709 = 1'b0;
    wire _707 = 1'b0;
    wire _706 = 1'b0;
    wire _704 = 1'b0;
    wire _703 = 1'b0;
    wire _701 = 1'b0;
    wire _700 = 1'b0;
    wire _698 = 1'b0;
    wire _697 = 1'b0;
    wire _695 = 1'b0;
    wire _694 = 1'b0;
    reg _696;
    reg _699;
    reg _702;
    reg _705;
    reg _708;
    reg _711;
    reg _714;
    reg _717;
    reg _720;
    wire _749;
    wire _750;
    wire write_enable_34;
    wire _755;
    wire [131:0] _762;
    wire [63:0] _763;
    wire _691 = 1'b0;
    wire _690 = 1'b0;
    wire _693;
    wire _23;
    reg PHASE_7;
    wire [63:0] _775;
    wire [11:0] address_35;
    wire write_enable_35;
    wire [11:0] address_36;
    wire _962;
    wire read_enable_29;
    wire _960;
    wire write_enable_36;
    wire _964;
    wire [131:0] _969;
    wire [63:0] _970;
    wire [11:0] _955 = 12'b000000000000;
    wire [11:0] address_37;
    wire _953;
    wire write_enable_37;
    wire [63:0] _878;
    wire [63:0] _877;
    wire [63:0] _879;
    wire [63:0] _875;
    wire [63:0] _874;
    wire [63:0] q1_2;
    wire [63:0] _880;
    wire [11:0] address_38;
    wire write_enable_38 = 1'b0;
    wire _865;
    wire read_enable_30;
    wire [11:0] address_39;
    wire _861;
    wire read_enable_31;
    wire _859;
    wire write_enable_39;
    wire _863;
    wire [131:0] _870;
    wire [63:0] _871;
    wire [63:0] data_35 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_36;
    wire [11:0] _853 = 12'b000000000000;
    wire _851;
    wire _850;
    wire _849;
    wire _848;
    wire _847;
    wire _846;
    wire _845;
    wire _844;
    wire _843;
    wire _842;
    wire _841;
    wire _840;
    wire [11:0] _852;
    wire [11:0] address_40;
    wire write_enable_40 = 1'b0;
    wire _837;
    wire read_enable_32;
    wire [63:0] data_37;
    wire [63:0] data_38;
    wire _834;
    wire _833;
    wire _832;
    wire _831;
    wire _830;
    wire _829;
    wire _828;
    wire _827;
    wire _826;
    wire _825;
    wire _824;
    wire _823;
    wire [11:0] _835;
    wire [11:0] address_41;
    wire _820;
    wire read_enable_33;
    wire _818;
    wire write_enable_41;
    wire _822;
    wire [131:0] _857;
    wire [63:0] _858;
    wire _777 = 1'b0;
    wire _776 = 1'b0;
    wire _779;
    wire _27;
    reg PHASE_8;
    wire [63:0] _872;
    wire [11:0] address_42;
    wire _810;
    wire read_enable_34;
    wire write_enable_42;
    wire _812;
    wire [11:0] address_43;
    wire _805;
    wire read_enable_35;
    wire _803;
    wire write_enable_43;
    wire _807;
    wire [131:0] _815;
    wire [63:0] _816;
    wire [63:0] _883;
    wire [63:0] data_39;
    wire [63:0] data_40;
    wire [63:0] data_41;
    wire [63:0] data_42;
    wire [11:0] address_44;
    wire _796;
    wire read_enable_36;
    wire _793;
    wire _794;
    wire write_enable_44;
    wire _798;
    wire [11:0] address_45;
    wire _789;
    wire read_enable_37;
    wire _786;
    wire _787;
    wire write_enable_45;
    wire _791;
    wire [131:0] _801;
    wire [63:0] _802;
    wire _784 = 1'b0;
    wire _783 = 1'b0;
    wire _884;
    wire _29;
    reg PHASE_9;
    wire [63:0] q0_2;
    wire _781 = 1'b0;
    wire _780 = 1'b0;
    reg _782;
    wire [63:0] _873;
    wire [191:0] _882;
    wire [63:0] _885;
    wire [63:0] data_43;
    wire [63:0] data_44;
    wire [63:0] data_45;
    wire [63:0] data_46;
    wire [11:0] address_46;
    wire _949;
    wire _948;
    wire read_enable_38;
    wire _942 = 1'b0;
    wire _941 = 1'b0;
    wire _939 = 1'b0;
    wire _938 = 1'b0;
    wire _936 = 1'b0;
    wire _935 = 1'b0;
    wire _933 = 1'b0;
    wire _932 = 1'b0;
    wire _930 = 1'b0;
    wire _929 = 1'b0;
    wire _927 = 1'b0;
    wire _926 = 1'b0;
    wire _924 = 1'b0;
    wire _923 = 1'b0;
    wire _921 = 1'b0;
    wire _920 = 1'b0;
    wire _918 = 1'b0;
    wire _917 = 1'b0;
    reg _919;
    reg _922;
    reg _925;
    reg _928;
    reg _931;
    reg _934;
    reg _937;
    reg _940;
    reg _943;
    wire _944;
    wire _915 = 1'b0;
    wire _914 = 1'b0;
    wire _912 = 1'b0;
    wire _911 = 1'b0;
    wire _909 = 1'b0;
    wire _908 = 1'b0;
    wire _906 = 1'b0;
    wire _905 = 1'b0;
    wire _903 = 1'b0;
    wire _902 = 1'b0;
    wire _900 = 1'b0;
    wire _899 = 1'b0;
    wire _897 = 1'b0;
    wire _896 = 1'b0;
    wire _894 = 1'b0;
    wire _893 = 1'b0;
    wire _891 = 1'b0;
    wire _890 = 1'b0;
    reg _892;
    reg _895;
    reg _898;
    reg _901;
    reg _904;
    reg _907;
    reg _910;
    reg _913;
    reg _916;
    wire _945;
    wire _946;
    wire write_enable_46;
    wire _951;
    wire [131:0] _958;
    wire [63:0] _959;
    wire _887 = 1'b0;
    wire _886 = 1'b0;
    wire _889;
    wire _31;
    reg PHASE_10;
    wire [63:0] _971;
    wire [11:0] address_47;
    wire write_enable_47;
    wire [11:0] address_48;
    wire _1158;
    wire read_enable_39;
    wire _1156;
    wire write_enable_48;
    wire _1160;
    wire [131:0] _1165;
    wire [63:0] _1166;
    wire [11:0] _1151 = 12'b000000000000;
    wire [11:0] address_49;
    wire _1149;
    wire write_enable_49;
    wire [63:0] _1074;
    wire [63:0] _1073;
    wire [63:0] _1075;
    wire [63:0] _1071;
    wire [63:0] _1070;
    wire [63:0] q1_3;
    wire [63:0] _1076;
    wire [11:0] address_50;
    wire write_enable_50 = 1'b0;
    wire _1061;
    wire read_enable_40;
    wire [11:0] address_51;
    wire _1057;
    wire read_enable_41;
    wire _1055;
    wire write_enable_51;
    wire _1059;
    wire [131:0] _1066;
    wire [63:0] _1067;
    wire [63:0] data_47 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_48;
    wire [11:0] _1049 = 12'b000000000000;
    wire _1047;
    wire _1046;
    wire _1045;
    wire _1044;
    wire _1043;
    wire _1042;
    wire _1041;
    wire _1040;
    wire _1039;
    wire _1038;
    wire _1037;
    wire _1036;
    wire [11:0] _1048;
    wire [11:0] address_52;
    wire write_enable_52 = 1'b0;
    wire _1033;
    wire read_enable_42;
    wire [63:0] data_49;
    wire [63:0] data_50;
    wire _1030;
    wire _1029;
    wire _1028;
    wire _1027;
    wire _1026;
    wire _1025;
    wire _1024;
    wire _1023;
    wire _1022;
    wire _1021;
    wire _1020;
    wire _1019;
    wire [11:0] _1031;
    wire [11:0] address_53;
    wire _1016;
    wire read_enable_43;
    wire _1014;
    wire write_enable_53;
    wire _1018;
    wire [131:0] _1053;
    wire [63:0] _1054;
    wire _973 = 1'b0;
    wire _972 = 1'b0;
    wire _975;
    wire _35;
    reg PHASE_11;
    wire [63:0] _1068;
    wire [11:0] address_54;
    wire _1006;
    wire read_enable_44;
    wire write_enable_54;
    wire _1008;
    wire [11:0] address_55;
    wire _1001;
    wire read_enable_45;
    wire _999;
    wire write_enable_55;
    wire _1003;
    wire [131:0] _1011;
    wire [63:0] _1012;
    wire [63:0] _1079;
    wire [63:0] data_51;
    wire [63:0] data_52;
    wire [63:0] data_53;
    wire [63:0] data_54;
    wire [11:0] address_56;
    wire _992;
    wire read_enable_46;
    wire _989;
    wire _990;
    wire write_enable_56;
    wire _994;
    wire [11:0] address_57;
    wire _985;
    wire read_enable_47;
    wire _982;
    wire _983;
    wire write_enable_57;
    wire _987;
    wire [131:0] _997;
    wire [63:0] _998;
    wire _980 = 1'b0;
    wire _979 = 1'b0;
    wire _1080;
    wire _37;
    reg PHASE_12;
    wire [63:0] q0_3;
    wire _977 = 1'b0;
    wire _976 = 1'b0;
    reg _978;
    wire [63:0] _1069;
    wire [191:0] _1078;
    wire [63:0] _1081;
    wire [63:0] data_55;
    wire [63:0] data_56;
    wire [63:0] data_57;
    wire [63:0] data_58;
    wire [11:0] address_58;
    wire _1145;
    wire _1144;
    wire read_enable_48;
    wire _1138 = 1'b0;
    wire _1137 = 1'b0;
    wire _1135 = 1'b0;
    wire _1134 = 1'b0;
    wire _1132 = 1'b0;
    wire _1131 = 1'b0;
    wire _1129 = 1'b0;
    wire _1128 = 1'b0;
    wire _1126 = 1'b0;
    wire _1125 = 1'b0;
    wire _1123 = 1'b0;
    wire _1122 = 1'b0;
    wire _1120 = 1'b0;
    wire _1119 = 1'b0;
    wire _1117 = 1'b0;
    wire _1116 = 1'b0;
    wire _1114 = 1'b0;
    wire _1113 = 1'b0;
    reg _1115;
    reg _1118;
    reg _1121;
    reg _1124;
    reg _1127;
    reg _1130;
    reg _1133;
    reg _1136;
    reg _1139;
    wire _1140;
    wire _1111 = 1'b0;
    wire _1110 = 1'b0;
    wire _1108 = 1'b0;
    wire _1107 = 1'b0;
    wire _1105 = 1'b0;
    wire _1104 = 1'b0;
    wire _1102 = 1'b0;
    wire _1101 = 1'b0;
    wire _1099 = 1'b0;
    wire _1098 = 1'b0;
    wire _1096 = 1'b0;
    wire _1095 = 1'b0;
    wire _1093 = 1'b0;
    wire _1092 = 1'b0;
    wire _1090 = 1'b0;
    wire _1089 = 1'b0;
    wire _1087 = 1'b0;
    wire _1086 = 1'b0;
    reg _1088;
    reg _1091;
    reg _1094;
    reg _1097;
    reg _1100;
    reg _1103;
    reg _1106;
    reg _1109;
    reg _1112;
    wire _1141;
    wire _1142;
    wire write_enable_58;
    wire _1147;
    wire [131:0] _1154;
    wire [63:0] _1155;
    wire _1083 = 1'b0;
    wire _1082 = 1'b0;
    wire _1085;
    wire _39;
    reg PHASE_13;
    wire [63:0] _1167;
    wire [11:0] address_59;
    wire write_enable_59;
    wire [11:0] address_60;
    wire _1354;
    wire read_enable_49;
    wire _1352;
    wire write_enable_60;
    wire _1356;
    wire [131:0] _1361;
    wire [63:0] _1362;
    wire [11:0] _1347 = 12'b000000000000;
    wire [11:0] address_61;
    wire _1345;
    wire write_enable_61;
    wire [63:0] _1270;
    wire [63:0] _1269;
    wire [63:0] _1271;
    wire [63:0] _1267;
    wire [63:0] _1266;
    wire [63:0] q1_4;
    wire [63:0] _1272;
    wire [11:0] address_62;
    wire write_enable_62 = 1'b0;
    wire _1257;
    wire read_enable_50;
    wire [11:0] address_63;
    wire _1253;
    wire read_enable_51;
    wire _1251;
    wire write_enable_63;
    wire _1255;
    wire [131:0] _1262;
    wire [63:0] _1263;
    wire [63:0] data_59 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_60;
    wire [11:0] _1245 = 12'b000000000000;
    wire _1243;
    wire _1242;
    wire _1241;
    wire _1240;
    wire _1239;
    wire _1238;
    wire _1237;
    wire _1236;
    wire _1235;
    wire _1234;
    wire _1233;
    wire _1232;
    wire [11:0] _1244;
    wire [11:0] address_64;
    wire write_enable_64 = 1'b0;
    wire _1229;
    wire read_enable_52;
    wire [63:0] data_61;
    wire [63:0] data_62;
    wire _1226;
    wire _1225;
    wire _1224;
    wire _1223;
    wire _1222;
    wire _1221;
    wire _1220;
    wire _1219;
    wire _1218;
    wire _1217;
    wire _1216;
    wire _1215;
    wire [11:0] _1227;
    wire [11:0] address_65;
    wire _1212;
    wire read_enable_53;
    wire _1210;
    wire write_enable_65;
    wire _1214;
    wire [131:0] _1249;
    wire [63:0] _1250;
    wire _1169 = 1'b0;
    wire _1168 = 1'b0;
    wire _1171;
    wire _43;
    reg PHASE_14;
    wire [63:0] _1264;
    wire [11:0] address_66;
    wire _1202;
    wire read_enable_54;
    wire write_enable_66;
    wire _1204;
    wire [11:0] address_67;
    wire _1197;
    wire read_enable_55;
    wire _1195;
    wire write_enable_67;
    wire _1199;
    wire [131:0] _1207;
    wire [63:0] _1208;
    wire [63:0] _1275;
    wire [63:0] data_63;
    wire [63:0] data_64;
    wire [63:0] data_65;
    wire [63:0] data_66;
    wire [11:0] address_68;
    wire _1188;
    wire read_enable_56;
    wire _1185;
    wire _1186;
    wire write_enable_68;
    wire _1190;
    wire [11:0] address_69;
    wire _1181;
    wire read_enable_57;
    wire _1178;
    wire _1179;
    wire write_enable_69;
    wire _1183;
    wire [131:0] _1193;
    wire [63:0] _1194;
    wire _1176 = 1'b0;
    wire _1175 = 1'b0;
    wire _1276;
    wire _45;
    reg PHASE_15;
    wire [63:0] q0_4;
    wire _1173 = 1'b0;
    wire _1172 = 1'b0;
    reg _1174;
    wire [63:0] _1265;
    wire [191:0] _1274;
    wire [63:0] _1277;
    wire [63:0] data_67;
    wire [63:0] data_68;
    wire [63:0] data_69;
    wire [63:0] data_70;
    wire [11:0] address_70;
    wire _1341;
    wire _1340;
    wire read_enable_58;
    wire _1334 = 1'b0;
    wire _1333 = 1'b0;
    wire _1331 = 1'b0;
    wire _1330 = 1'b0;
    wire _1328 = 1'b0;
    wire _1327 = 1'b0;
    wire _1325 = 1'b0;
    wire _1324 = 1'b0;
    wire _1322 = 1'b0;
    wire _1321 = 1'b0;
    wire _1319 = 1'b0;
    wire _1318 = 1'b0;
    wire _1316 = 1'b0;
    wire _1315 = 1'b0;
    wire _1313 = 1'b0;
    wire _1312 = 1'b0;
    wire _1310 = 1'b0;
    wire _1309 = 1'b0;
    reg _1311;
    reg _1314;
    reg _1317;
    reg _1320;
    reg _1323;
    reg _1326;
    reg _1329;
    reg _1332;
    reg _1335;
    wire _1336;
    wire _1307 = 1'b0;
    wire _1306 = 1'b0;
    wire _1304 = 1'b0;
    wire _1303 = 1'b0;
    wire _1301 = 1'b0;
    wire _1300 = 1'b0;
    wire _1298 = 1'b0;
    wire _1297 = 1'b0;
    wire _1295 = 1'b0;
    wire _1294 = 1'b0;
    wire _1292 = 1'b0;
    wire _1291 = 1'b0;
    wire _1289 = 1'b0;
    wire _1288 = 1'b0;
    wire _1286 = 1'b0;
    wire _1285 = 1'b0;
    wire _1283 = 1'b0;
    wire _1282 = 1'b0;
    reg _1284;
    reg _1287;
    reg _1290;
    reg _1293;
    reg _1296;
    reg _1299;
    reg _1302;
    reg _1305;
    reg _1308;
    wire _1337;
    wire _1338;
    wire write_enable_70;
    wire _1343;
    wire [131:0] _1350;
    wire [63:0] _1351;
    wire _1279 = 1'b0;
    wire _1278 = 1'b0;
    wire _1281;
    wire _47;
    reg PHASE_16;
    wire [63:0] _1363;
    wire [11:0] address_71;
    wire write_enable_71;
    wire [11:0] address_72;
    wire _1550;
    wire read_enable_59;
    wire _1548;
    wire write_enable_72;
    wire _1552;
    wire [131:0] _1557;
    wire [63:0] _1558;
    wire [11:0] _1543 = 12'b000000000000;
    wire [11:0] address_73;
    wire _1541;
    wire write_enable_73;
    wire [63:0] _1466;
    wire [63:0] _1465;
    wire [63:0] _1467;
    wire [63:0] _1463;
    wire [63:0] _1462;
    wire [63:0] q1_5;
    wire [63:0] _1468;
    wire [11:0] address_74;
    wire write_enable_74 = 1'b0;
    wire _1453;
    wire read_enable_60;
    wire [11:0] address_75;
    wire _1449;
    wire read_enable_61;
    wire _1447;
    wire write_enable_75;
    wire _1451;
    wire [131:0] _1458;
    wire [63:0] _1459;
    wire [63:0] data_71 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_72;
    wire [11:0] _1441 = 12'b000000000000;
    wire _1439;
    wire _1438;
    wire _1437;
    wire _1436;
    wire _1435;
    wire _1434;
    wire _1433;
    wire _1432;
    wire _1431;
    wire _1430;
    wire _1429;
    wire _1428;
    wire [11:0] _1440;
    wire [11:0] address_76;
    wire write_enable_76 = 1'b0;
    wire _1425;
    wire read_enable_62;
    wire [63:0] data_73;
    wire [63:0] data_74;
    wire _1422;
    wire _1421;
    wire _1420;
    wire _1419;
    wire _1418;
    wire _1417;
    wire _1416;
    wire _1415;
    wire _1414;
    wire _1413;
    wire _1412;
    wire _1411;
    wire [11:0] _1423;
    wire [11:0] address_77;
    wire _1408;
    wire read_enable_63;
    wire _1406;
    wire write_enable_77;
    wire _1410;
    wire [131:0] _1445;
    wire [63:0] _1446;
    wire _1365 = 1'b0;
    wire _1364 = 1'b0;
    wire _1367;
    wire _51;
    reg PHASE_17;
    wire [63:0] _1460;
    wire [11:0] address_78;
    wire _1398;
    wire read_enable_64;
    wire write_enable_78;
    wire _1400;
    wire [11:0] address_79;
    wire _1393;
    wire read_enable_65;
    wire _1391;
    wire write_enable_79;
    wire _1395;
    wire [131:0] _1403;
    wire [63:0] _1404;
    wire [63:0] _1471;
    wire [63:0] data_75;
    wire [63:0] data_76;
    wire [63:0] data_77;
    wire [63:0] data_78;
    wire [11:0] address_80;
    wire _1384;
    wire read_enable_66;
    wire _1381;
    wire _1382;
    wire write_enable_80;
    wire _1386;
    wire [11:0] address_81;
    wire _1377;
    wire read_enable_67;
    wire _1374;
    wire _1375;
    wire write_enable_81;
    wire _1379;
    wire [131:0] _1389;
    wire [63:0] _1390;
    wire _1372 = 1'b0;
    wire _1371 = 1'b0;
    wire _1472;
    wire _53;
    reg PHASE_18;
    wire [63:0] q0_5;
    wire _1369 = 1'b0;
    wire _1368 = 1'b0;
    reg _1370;
    wire [63:0] _1461;
    wire [191:0] _1470;
    wire [63:0] _1473;
    wire [63:0] data_79;
    wire [63:0] data_80;
    wire [63:0] data_81;
    wire [63:0] data_82;
    wire [11:0] address_82;
    wire _1537;
    wire _1536;
    wire read_enable_68;
    wire _1530 = 1'b0;
    wire _1529 = 1'b0;
    wire _1527 = 1'b0;
    wire _1526 = 1'b0;
    wire _1524 = 1'b0;
    wire _1523 = 1'b0;
    wire _1521 = 1'b0;
    wire _1520 = 1'b0;
    wire _1518 = 1'b0;
    wire _1517 = 1'b0;
    wire _1515 = 1'b0;
    wire _1514 = 1'b0;
    wire _1512 = 1'b0;
    wire _1511 = 1'b0;
    wire _1509 = 1'b0;
    wire _1508 = 1'b0;
    wire _1506 = 1'b0;
    wire _1505 = 1'b0;
    reg _1507;
    reg _1510;
    reg _1513;
    reg _1516;
    reg _1519;
    reg _1522;
    reg _1525;
    reg _1528;
    reg _1531;
    wire _1532;
    wire _1503 = 1'b0;
    wire _1502 = 1'b0;
    wire _1500 = 1'b0;
    wire _1499 = 1'b0;
    wire _1497 = 1'b0;
    wire _1496 = 1'b0;
    wire _1494 = 1'b0;
    wire _1493 = 1'b0;
    wire _1491 = 1'b0;
    wire _1490 = 1'b0;
    wire _1488 = 1'b0;
    wire _1487 = 1'b0;
    wire _1485 = 1'b0;
    wire _1484 = 1'b0;
    wire _1482 = 1'b0;
    wire _1481 = 1'b0;
    wire _1479 = 1'b0;
    wire _1478 = 1'b0;
    reg _1480;
    reg _1483;
    reg _1486;
    reg _1489;
    reg _1492;
    reg _1495;
    reg _1498;
    reg _1501;
    reg _1504;
    wire _1533;
    wire _1534;
    wire write_enable_82;
    wire _1539;
    wire [131:0] _1546;
    wire [63:0] _1547;
    wire _1475 = 1'b0;
    wire _1474 = 1'b0;
    wire _1477;
    wire _55;
    reg PHASE_19;
    wire [63:0] _1559;
    wire [11:0] address_83;
    wire write_enable_83;
    wire [11:0] address_84;
    wire _1746;
    wire read_enable_69;
    wire _1744;
    wire write_enable_84;
    wire _1748;
    wire [131:0] _1753;
    wire [63:0] _1754;
    wire [11:0] _1739 = 12'b000000000000;
    wire [11:0] address_85;
    wire _1737;
    wire write_enable_85;
    wire [3:0] _292;
    wire _291;
    wire _289;
    wire [63:0] _288;
    wire [63:0] _287;
    wire [63:0] _286;
    wire [63:0] _285;
    wire [63:0] _284;
    wire [63:0] _283;
    wire [63:0] _282;
    wire [63:0] _1662;
    wire [63:0] _1661;
    wire [63:0] _1663;
    wire [63:0] _1659;
    wire [63:0] _1658;
    wire [63:0] q1_6;
    wire [63:0] _1664;
    wire [11:0] address_86;
    wire write_enable_86 = 1'b0;
    wire _1649;
    wire read_enable_70;
    wire [11:0] address_87;
    wire _1645;
    wire read_enable_71;
    wire _1643;
    wire write_enable_87;
    wire _1647;
    wire [131:0] _1654;
    wire [63:0] _1655;
    wire [63:0] data_83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_84;
    wire [11:0] _1637 = 12'b000000000000;
    wire _1635;
    wire _1634;
    wire _1633;
    wire _1632;
    wire _1631;
    wire _1630;
    wire _1629;
    wire _1628;
    wire _1627;
    wire _1626;
    wire _1625;
    wire _1624;
    wire [11:0] _1636;
    wire [11:0] address_88;
    wire write_enable_88 = 1'b0;
    wire _1621;
    wire read_enable_72;
    wire [63:0] data_85;
    wire [63:0] data_86;
    wire [11:0] _60;
    wire _1618;
    wire _1617;
    wire _1616;
    wire _1615;
    wire _1614;
    wire _1613;
    wire _1612;
    wire _1611;
    wire _1610;
    wire _1609;
    wire _1608;
    wire _1607;
    wire [11:0] _1619;
    wire [11:0] address_89;
    wire _1604;
    wire read_enable_73;
    wire [7:0] _62;
    wire _1602;
    wire write_enable_89;
    wire _1606;
    wire [131:0] _1641;
    wire [63:0] _1642;
    wire _1561 = 1'b0;
    wire _1560 = 1'b0;
    wire _1563;
    wire _63;
    reg PHASE_20;
    wire [63:0] _1656;
    wire [11:0] address_90;
    wire _1594;
    wire read_enable_74;
    wire write_enable_90;
    wire _1596;
    wire [11:0] address_91;
    wire _1589;
    wire read_enable_75;
    wire _1587;
    wire write_enable_91;
    wire _1591;
    wire [131:0] _1599;
    wire [63:0] _1600;
    wire [63:0] _1667;
    wire [63:0] data_87;
    wire [63:0] data_88;
    wire [63:0] data_89;
    wire [63:0] data_90;
    wire [11:0] _198 = 12'b000000000000;
    wire [11:0] _197 = 12'b000000000000;
    wire [11:0] _195 = 12'b000000000000;
    wire [11:0] _194 = 12'b000000000000;
    wire [11:0] _192 = 12'b000000000000;
    wire [11:0] _191 = 12'b000000000000;
    wire [11:0] _189 = 12'b000000000000;
    wire [11:0] _188 = 12'b000000000000;
    wire [11:0] _186 = 12'b000000000000;
    wire [11:0] _185 = 12'b000000000000;
    wire [11:0] _183 = 12'b000000000000;
    wire [11:0] _182 = 12'b000000000000;
    wire [11:0] _180 = 12'b000000000000;
    wire [11:0] _179 = 12'b000000000000;
    wire [11:0] _177 = 12'b000000000000;
    wire [11:0] _176 = 12'b000000000000;
    wire [11:0] _174 = 12'b000000000000;
    wire [11:0] _173 = 12'b000000000000;
    reg [11:0] _175;
    reg [11:0] _178;
    reg [11:0] _181;
    reg [11:0] _184;
    reg [11:0] _187;
    reg [11:0] _190;
    reg [11:0] _193;
    reg [11:0] _196;
    reg [11:0] _199;
    wire [11:0] _172;
    wire [11:0] address_92;
    wire _1580;
    wire read_enable_76;
    wire _1577;
    wire _1578;
    wire write_enable_92;
    wire _1582;
    wire [11:0] address_93;
    wire _1573;
    wire read_enable_77;
    wire _1570;
    wire _1571;
    wire write_enable_93;
    wire _1575;
    wire [131:0] _1585;
    wire [63:0] _1586;
    wire _99;
    wire _1568 = 1'b0;
    wire _1567 = 1'b0;
    wire _1668;
    wire _65;
    reg PHASE_21;
    wire [63:0] q0_6;
    wire _1565 = 1'b0;
    wire _1564 = 1'b0;
    wire _92;
    reg _1566;
    wire [63:0] _1657;
    wire [191:0] _1666;
    wire [63:0] _1669;
    wire [63:0] data_91;
    wire [63:0] data_92;
    wire [63:0] data_93;
    wire [63:0] data_94;
    wire [11:0] _163 = 12'b000000000000;
    wire [11:0] _162 = 12'b000000000000;
    wire [11:0] _160 = 12'b000000000000;
    wire [11:0] _159 = 12'b000000000000;
    wire [11:0] _157 = 12'b000000000000;
    wire [11:0] _156 = 12'b000000000000;
    wire [11:0] _154 = 12'b000000000000;
    wire [11:0] _153 = 12'b000000000000;
    wire [11:0] _151 = 12'b000000000000;
    wire [11:0] _150 = 12'b000000000000;
    wire [11:0] _148 = 12'b000000000000;
    wire [11:0] _147 = 12'b000000000000;
    wire [11:0] _145 = 12'b000000000000;
    wire [11:0] _144 = 12'b000000000000;
    wire [11:0] _142 = 12'b000000000000;
    wire [11:0] _141 = 12'b000000000000;
    wire [11:0] _139 = 12'b000000000000;
    wire [11:0] _138 = 12'b000000000000;
    wire [11:0] _137;
    reg [11:0] _140;
    reg [11:0] _143;
    reg [11:0] _146;
    reg [11:0] _149;
    reg [11:0] _152;
    reg [11:0] _155;
    reg [11:0] _158;
    reg [11:0] _161;
    reg [11:0] _164;
    wire [11:0] _68;
    wire [11:0] address_94;
    wire _1733;
    wire [7:0] _70;
    wire _1732;
    wire read_enable_78;
    wire _1726 = 1'b0;
    wire _1725 = 1'b0;
    wire _1723 = 1'b0;
    wire _1722 = 1'b0;
    wire _1720 = 1'b0;
    wire _1719 = 1'b0;
    wire _1717 = 1'b0;
    wire _1716 = 1'b0;
    wire _1714 = 1'b0;
    wire _1713 = 1'b0;
    wire _1711 = 1'b0;
    wire _1710 = 1'b0;
    wire _1708 = 1'b0;
    wire _1707 = 1'b0;
    wire _1705 = 1'b0;
    wire _1704 = 1'b0;
    wire _1702 = 1'b0;
    wire _1701 = 1'b0;
    wire _290;
    reg _1703;
    reg _1706;
    reg _1709;
    reg _1712;
    reg _1715;
    reg _1718;
    reg _1721;
    reg _1724;
    reg _1727;
    wire _1728;
    wire _1699 = 1'b0;
    wire _1698 = 1'b0;
    wire _1696 = 1'b0;
    wire _1695 = 1'b0;
    wire _1693 = 1'b0;
    wire _1692 = 1'b0;
    wire _1690 = 1'b0;
    wire _1689 = 1'b0;
    wire _1687 = 1'b0;
    wire _1686 = 1'b0;
    wire _1684 = 1'b0;
    wire _1683 = 1'b0;
    wire _1681 = 1'b0;
    wire _1680 = 1'b0;
    wire _1678 = 1'b0;
    wire _1677 = 1'b0;
    wire _1675 = 1'b0;
    wire _1674 = 1'b0;
    wire _130;
    reg _1676;
    reg _1679;
    reg _1682;
    reg _1685;
    reg _1688;
    reg _1691;
    reg _1694;
    reg _1697;
    reg _1700;
    wire _1729;
    wire _128 = 1'b0;
    wire _127 = 1'b0;
    wire _125 = 1'b0;
    wire _124 = 1'b0;
    wire _122 = 1'b0;
    wire _121 = 1'b0;
    wire _119 = 1'b0;
    wire _118 = 1'b0;
    wire _116 = 1'b0;
    wire _115 = 1'b0;
    wire _113 = 1'b0;
    wire _112 = 1'b0;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire vdd = 1'b1;
    wire _104 = 1'b0;
    wire _103 = 1'b0;
    wire _102;
    reg _105;
    reg _108;
    reg _111;
    reg _114;
    reg _117;
    reg _120;
    reg _123;
    reg _126;
    reg _129;
    wire _1730;
    wire write_enable_94;
    wire _1735;
    wire gnd = 1'b0;
    wire [131:0] _1742;
    wire [63:0] _1743;
    wire _72;
    wire _1671 = 1'b0;
    wire _1670 = 1'b0;
    wire _1673;
    wire _73;
    reg PHASE_22;
    wire [63:0] _1755;
    wire _76;
    wire _78;
    wire _80;
    wire _82;
    wire _84;
    wire [523:0] _91;
    wire _1756;

    /* logic */
    assign address = _372 ? _199 : _367;
    assign write_enable = _365 & _372;
    assign address_0 = _372 ? _164 : _68;
    assign _374 = ~ _372;
    assign read_enable = _360 & _374;
    assign _372 = ~ PHASE_1;
    assign write_enable_0 = _358 & _372;
    assign _376 = write_enable_0 | read_enable;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_376), .regcea(vdd), .wea(write_enable_0), .addra(address_0), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable), .regceb(vdd), .web(write_enable), .addrb(address), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_381[131:131]), .sbiterrb(_381[130:130]), .doutb(_381[129:66]), .dbiterra(_381[65:65]), .sbiterra(_381[64:64]), .douta(_381[63:0]) );
    assign _382 = _381[63:0];
    assign address_1 = PHASE_1 ? _199 : _367;
    assign _365 = _129 & _328;
    assign write_enable_1 = _365 & PHASE_1;
    assign _279 = _271[129:66];
    assign _278 = _258[129:66];
    assign _280 = PHASE ? _279 : _278;
    assign _276 = _216[129:66];
    assign _275 = _202[129:66];
    assign q1 = PHASE_0 ? _276 : _275;
    assign _281 = _96 ? _280 : q1;
    assign address_2 = _260 ? _254 : _253;
    assign _266 = ~ _260;
    assign read_enable_0 = _102 & _266;
    assign address_3 = _260 ? _60 : _236;
    assign _262 = ~ _260;
    assign read_enable_1 = _102 & _262;
    assign _260 = ~ PHASE;
    assign write_enable_3 = _219 & _260;
    assign _264 = write_enable_3 | read_enable_1;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_0
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_264), .regcea(vdd), .wea(write_enable_3), .addra(address_3), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_0), .regceb(vdd), .web(write_enable_2), .addrb(address_2), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_271[131:131]), .sbiterrb(_271[130:130]), .doutb(_271[129:66]), .dbiterra(_271[65:65]), .sbiterra(_271[64:64]), .douta(_271[63:0]) );
    assign _272 = _271[63:0];
    assign _252 = _172[11:11];
    assign _251 = _172[10:10];
    assign _250 = _172[9:9];
    assign _249 = _172[8:8];
    assign _248 = _172[7:7];
    assign _247 = _172[6:6];
    assign _246 = _172[5:5];
    assign _245 = _172[4:4];
    assign _244 = _172[3:3];
    assign _243 = _172[2:2];
    assign _242 = _172[1:1];
    assign _241 = _172[0:0];
    assign _253 = { _241, _242, _243, _244, _245, _246, _247, _248, _249, _250, _251, _252 };
    assign address_4 = PHASE ? _254 : _253;
    assign _238 = ~ PHASE;
    assign read_enable_2 = _102 & _238;
    assign data_1 = wr_d7;
    assign _235 = _137[11:11];
    assign _234 = _137[10:10];
    assign _233 = _137[9:9];
    assign _232 = _137[8:8];
    assign _231 = _137[7:7];
    assign _230 = _137[6:6];
    assign _229 = _137[5:5];
    assign _228 = _137[4:4];
    assign _227 = _137[3:3];
    assign _226 = _137[2:2];
    assign _225 = _137[1:1];
    assign _224 = _137[0:0];
    assign _236 = { _224, _225, _226, _227, _228, _229, _230, _231, _232, _233, _234, _235 };
    assign address_5 = PHASE ? _60 : _236;
    assign _221 = ~ PHASE;
    assign read_enable_3 = _102 & _221;
    assign _219 = _62[7:7];
    assign write_enable_5 = _219 & PHASE;
    assign _223 = write_enable_5 | read_enable_3;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_1
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_223), .regcea(vdd), .wea(write_enable_5), .addra(address_5), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_2), .regceb(vdd), .web(write_enable_4), .addrb(address_4), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_258[131:131]), .sbiterrb(_258[130:130]), .doutb(_258[129:66]), .dbiterra(_258[65:65]), .sbiterra(_258[64:64]), .douta(_258[63:0]) );
    assign _259 = _258[63:0];
    assign _89 = ~ PHASE;
    assign _3 = _89;
    always @(posedge _84) begin
        if (_82)
            PHASE <= _87;
        else
            if (_72)
                PHASE <= _3;
    end
    assign _273 = PHASE ? _272 : _259;
    assign address_6 = _204 ? _199 : _172;
    assign _211 = ~ _204;
    assign read_enable_4 = _102 & _211;
    assign write_enable_6 = _167 & _204;
    assign _213 = write_enable_6 | read_enable_4;
    assign address_7 = _204 ? _164 : _137;
    assign _206 = ~ _204;
    assign read_enable_5 = _102 & _206;
    assign _204 = ~ PHASE_0;
    assign write_enable_7 = _132 & _204;
    assign _208 = write_enable_7 | read_enable_5;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_2
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_208), .regcea(vdd), .wea(write_enable_7), .addra(address_7), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_213), .regceb(vdd), .web(write_enable_6), .addrb(address_6), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_216[131:131]), .sbiterrb(_216[130:130]), .doutb(_216[129:66]), .dbiterra(_216[65:65]), .sbiterra(_216[64:64]), .douta(_216[63:0]) );
    assign _217 = _216[63:0];
    assign _295 = _294[127:64];
    assign data_3 = _295;
    assign address_8 = PHASE_0 ? _199 : _172;
    assign _169 = ~ PHASE_0;
    assign read_enable_6 = _102 & _169;
    assign _166 = ~ _130;
    assign _167 = _129 & _166;
    assign write_enable_8 = _167 & PHASE_0;
    assign _171 = write_enable_8 | read_enable_6;
    assign address_9 = PHASE_0 ? _164 : _137;
    assign _134 = ~ PHASE_0;
    assign read_enable_7 = _102 & _134;
    assign _131 = ~ _130;
    assign _132 = _129 & _131;
    assign write_enable_9 = _132 & PHASE_0;
    assign _136 = write_enable_9 | read_enable_7;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_3
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_136), .regcea(vdd), .wea(write_enable_9), .addra(address_9), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_171), .regceb(vdd), .web(write_enable_8), .addrb(address_8), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_202[131:131]), .sbiterrb(_202[130:130]), .doutb(_202[129:66]), .dbiterra(_202[65:65]), .sbiterra(_202[64:64]), .douta(_202[63:0]) );
    assign _203 = _202[63:0];
    assign _296 = ~ PHASE_0;
    assign _5 = _296;
    always @(posedge _84) begin
        if (_82)
            PHASE_0 <= _98;
        else
            if (_99)
                PHASE_0 <= _5;
    end
    assign q0 = PHASE_0 ? _217 : _203;
    always @(posedge _84) begin
        if (_82)
            _96 <= _94;
        else
            _96 <= _92;
    end
    assign _274 = _96 ? _273 : q0;
    dp_38
        dp_6
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_274), .d2(_281), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_294[191:128]), .q2(_294[127:64]), .q1(_294[63:0]) );
    assign _297 = _294[63:0];
    assign data_7 = _297;
    assign address_10 = PHASE_1 ? _164 : _68;
    assign _361 = ~ PHASE_1;
    assign _360 = _70[7:7];
    assign read_enable_8 = _360 & _361;
    always @(posedge _84) begin
        if (_82)
            _331 <= _330;
        else
            _331 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _334 <= _333;
        else
            _334 <= _331;
    end
    always @(posedge _84) begin
        if (_82)
            _337 <= _336;
        else
            _337 <= _334;
    end
    always @(posedge _84) begin
        if (_82)
            _340 <= _339;
        else
            _340 <= _337;
    end
    always @(posedge _84) begin
        if (_82)
            _343 <= _342;
        else
            _343 <= _340;
    end
    always @(posedge _84) begin
        if (_82)
            _346 <= _345;
        else
            _346 <= _343;
    end
    always @(posedge _84) begin
        if (_82)
            _349 <= _348;
        else
            _349 <= _346;
    end
    always @(posedge _84) begin
        if (_82)
            _352 <= _351;
        else
            _352 <= _349;
    end
    always @(posedge _84) begin
        if (_82)
            _355 <= _354;
        else
            _355 <= _352;
    end
    assign _356 = ~ _355;
    always @(posedge _84) begin
        if (_82)
            _304 <= _303;
        else
            _304 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _307 <= _306;
        else
            _307 <= _304;
    end
    always @(posedge _84) begin
        if (_82)
            _310 <= _309;
        else
            _310 <= _307;
    end
    always @(posedge _84) begin
        if (_82)
            _313 <= _312;
        else
            _313 <= _310;
    end
    always @(posedge _84) begin
        if (_82)
            _316 <= _315;
        else
            _316 <= _313;
    end
    always @(posedge _84) begin
        if (_82)
            _319 <= _318;
        else
            _319 <= _316;
    end
    always @(posedge _84) begin
        if (_82)
            _322 <= _321;
        else
            _322 <= _319;
    end
    always @(posedge _84) begin
        if (_82)
            _325 <= _324;
        else
            _325 <= _322;
    end
    always @(posedge _84) begin
        if (_82)
            _328 <= _327;
        else
            _328 <= _325;
    end
    assign _357 = _328 & _356;
    assign _358 = _129 & _357;
    assign write_enable_10 = _358 & PHASE_1;
    assign _363 = write_enable_10 | read_enable_8;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_4
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_363), .regcea(vdd), .wea(write_enable_10), .addra(address_10), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_1), .regceb(vdd), .web(write_enable_1), .addrb(address_1), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_370[131:131]), .sbiterrb(_370[130:130]), .doutb(_370[129:66]), .dbiterra(_370[65:65]), .sbiterra(_370[64:64]), .douta(_370[63:0]) );
    assign _371 = _370[63:0];
    assign _301 = ~ PHASE_1;
    assign _7 = _301;
    always @(posedge _84) begin
        if (_82)
            PHASE_1 <= _299;
        else
            if (_72)
                PHASE_1 <= _7;
    end
    assign _383 = PHASE_1 ? _382 : _371;
    assign address_11 = _568 ? _199 : _563;
    assign write_enable_11 = _561 & _568;
    assign address_12 = _568 ? _164 : _68;
    assign _570 = ~ _568;
    assign read_enable_9 = _556 & _570;
    assign _568 = ~ PHASE_4;
    assign write_enable_12 = _554 & _568;
    assign _572 = write_enable_12 | read_enable_9;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_5
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_572), .regcea(vdd), .wea(write_enable_12), .addra(address_12), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_11), .regceb(vdd), .web(write_enable_11), .addrb(address_11), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_577[131:131]), .sbiterrb(_577[130:130]), .doutb(_577[129:66]), .dbiterra(_577[65:65]), .sbiterra(_577[64:64]), .douta(_577[63:0]) );
    assign _578 = _577[63:0];
    assign address_13 = PHASE_4 ? _199 : _563;
    assign _561 = _129 & _524;
    assign write_enable_13 = _561 & PHASE_4;
    assign _486 = _478[129:66];
    assign _485 = _465[129:66];
    assign _487 = PHASE_2 ? _486 : _485;
    assign _483 = _423[129:66];
    assign _482 = _409[129:66];
    assign q1_0 = PHASE_3 ? _483 : _482;
    assign _488 = _390 ? _487 : q1_0;
    assign address_14 = _467 ? _461 : _460;
    assign _473 = ~ _467;
    assign read_enable_10 = _102 & _473;
    assign address_15 = _467 ? _60 : _443;
    assign _469 = ~ _467;
    assign read_enable_11 = _102 & _469;
    assign _467 = ~ PHASE_2;
    assign write_enable_15 = _426 & _467;
    assign _471 = write_enable_15 | read_enable_11;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_6
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_471), .regcea(vdd), .wea(write_enable_15), .addra(address_15), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_10), .regceb(vdd), .web(write_enable_14), .addrb(address_14), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_478[131:131]), .sbiterrb(_478[130:130]), .doutb(_478[129:66]), .dbiterra(_478[65:65]), .sbiterra(_478[64:64]), .douta(_478[63:0]) );
    assign _479 = _478[63:0];
    assign _459 = _172[11:11];
    assign _458 = _172[10:10];
    assign _457 = _172[9:9];
    assign _456 = _172[8:8];
    assign _455 = _172[7:7];
    assign _454 = _172[6:6];
    assign _453 = _172[5:5];
    assign _452 = _172[4:4];
    assign _451 = _172[3:3];
    assign _450 = _172[2:2];
    assign _449 = _172[1:1];
    assign _448 = _172[0:0];
    assign _460 = { _448, _449, _450, _451, _452, _453, _454, _455, _456, _457, _458, _459 };
    assign address_16 = PHASE_2 ? _461 : _460;
    assign _445 = ~ PHASE_2;
    assign read_enable_12 = _102 & _445;
    assign data_13 = wr_d6;
    assign _442 = _137[11:11];
    assign _441 = _137[10:10];
    assign _440 = _137[9:9];
    assign _439 = _137[8:8];
    assign _438 = _137[7:7];
    assign _437 = _137[6:6];
    assign _436 = _137[5:5];
    assign _435 = _137[4:4];
    assign _434 = _137[3:3];
    assign _433 = _137[2:2];
    assign _432 = _137[1:1];
    assign _431 = _137[0:0];
    assign _443 = { _431, _432, _433, _434, _435, _436, _437, _438, _439, _440, _441, _442 };
    assign address_17 = PHASE_2 ? _60 : _443;
    assign _428 = ~ PHASE_2;
    assign read_enable_13 = _102 & _428;
    assign _426 = _62[6:6];
    assign write_enable_17 = _426 & PHASE_2;
    assign _430 = write_enable_17 | read_enable_13;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_7
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_430), .regcea(vdd), .wea(write_enable_17), .addra(address_17), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_12), .regceb(vdd), .web(write_enable_16), .addrb(address_16), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_465[131:131]), .sbiterrb(_465[130:130]), .doutb(_465[129:66]), .dbiterra(_465[65:65]), .sbiterra(_465[64:64]), .douta(_465[63:0]) );
    assign _466 = _465[63:0];
    assign _387 = ~ PHASE_2;
    assign _11 = _387;
    always @(posedge _84) begin
        if (_82)
            PHASE_2 <= _385;
        else
            if (_72)
                PHASE_2 <= _11;
    end
    assign _480 = PHASE_2 ? _479 : _466;
    assign address_18 = _411 ? _199 : _172;
    assign _418 = ~ _411;
    assign read_enable_14 = _102 & _418;
    assign write_enable_18 = _402 & _411;
    assign _420 = write_enable_18 | read_enable_14;
    assign address_19 = _411 ? _164 : _137;
    assign _413 = ~ _411;
    assign read_enable_15 = _102 & _413;
    assign _411 = ~ PHASE_3;
    assign write_enable_19 = _395 & _411;
    assign _415 = write_enable_19 | read_enable_15;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_8
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_415), .regcea(vdd), .wea(write_enable_19), .addra(address_19), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_420), .regceb(vdd), .web(write_enable_18), .addrb(address_18), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_423[131:131]), .sbiterrb(_423[130:130]), .doutb(_423[129:66]), .dbiterra(_423[65:65]), .sbiterra(_423[64:64]), .douta(_423[63:0]) );
    assign _424 = _423[63:0];
    assign _491 = _490[127:64];
    assign data_15 = _491;
    assign address_20 = PHASE_3 ? _199 : _172;
    assign _404 = ~ PHASE_3;
    assign read_enable_16 = _102 & _404;
    assign _401 = ~ _130;
    assign _402 = _129 & _401;
    assign write_enable_20 = _402 & PHASE_3;
    assign _406 = write_enable_20 | read_enable_16;
    assign address_21 = PHASE_3 ? _164 : _137;
    assign _397 = ~ PHASE_3;
    assign read_enable_17 = _102 & _397;
    assign _394 = ~ _130;
    assign _395 = _129 & _394;
    assign write_enable_21 = _395 & PHASE_3;
    assign _399 = write_enable_21 | read_enable_17;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_9
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_399), .regcea(vdd), .wea(write_enable_21), .addra(address_21), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_406), .regceb(vdd), .web(write_enable_20), .addrb(address_20), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_409[131:131]), .sbiterrb(_409[130:130]), .doutb(_409[129:66]), .dbiterra(_409[65:65]), .sbiterra(_409[64:64]), .douta(_409[63:0]) );
    assign _410 = _409[63:0];
    assign _492 = ~ PHASE_3;
    assign _13 = _492;
    always @(posedge _84) begin
        if (_82)
            PHASE_3 <= _392;
        else
            if (_99)
                PHASE_3 <= _13;
    end
    assign q0_0 = PHASE_3 ? _424 : _410;
    always @(posedge _84) begin
        if (_82)
            _390 <= _389;
        else
            _390 <= _92;
    end
    assign _481 = _390 ? _480 : q0_0;
    dp_37
        dp_5
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_481), .d2(_488), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_490[191:128]), .q2(_490[127:64]), .q1(_490[63:0]) );
    assign _493 = _490[63:0];
    assign data_19 = _493;
    assign address_22 = PHASE_4 ? _164 : _68;
    assign _557 = ~ PHASE_4;
    assign _556 = _70[6:6];
    assign read_enable_18 = _556 & _557;
    always @(posedge _84) begin
        if (_82)
            _527 <= _526;
        else
            _527 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _530 <= _529;
        else
            _530 <= _527;
    end
    always @(posedge _84) begin
        if (_82)
            _533 <= _532;
        else
            _533 <= _530;
    end
    always @(posedge _84) begin
        if (_82)
            _536 <= _535;
        else
            _536 <= _533;
    end
    always @(posedge _84) begin
        if (_82)
            _539 <= _538;
        else
            _539 <= _536;
    end
    always @(posedge _84) begin
        if (_82)
            _542 <= _541;
        else
            _542 <= _539;
    end
    always @(posedge _84) begin
        if (_82)
            _545 <= _544;
        else
            _545 <= _542;
    end
    always @(posedge _84) begin
        if (_82)
            _548 <= _547;
        else
            _548 <= _545;
    end
    always @(posedge _84) begin
        if (_82)
            _551 <= _550;
        else
            _551 <= _548;
    end
    assign _552 = ~ _551;
    always @(posedge _84) begin
        if (_82)
            _500 <= _499;
        else
            _500 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _503 <= _502;
        else
            _503 <= _500;
    end
    always @(posedge _84) begin
        if (_82)
            _506 <= _505;
        else
            _506 <= _503;
    end
    always @(posedge _84) begin
        if (_82)
            _509 <= _508;
        else
            _509 <= _506;
    end
    always @(posedge _84) begin
        if (_82)
            _512 <= _511;
        else
            _512 <= _509;
    end
    always @(posedge _84) begin
        if (_82)
            _515 <= _514;
        else
            _515 <= _512;
    end
    always @(posedge _84) begin
        if (_82)
            _518 <= _517;
        else
            _518 <= _515;
    end
    always @(posedge _84) begin
        if (_82)
            _521 <= _520;
        else
            _521 <= _518;
    end
    always @(posedge _84) begin
        if (_82)
            _524 <= _523;
        else
            _524 <= _521;
    end
    assign _553 = _524 & _552;
    assign _554 = _129 & _553;
    assign write_enable_22 = _554 & PHASE_4;
    assign _559 = write_enable_22 | read_enable_18;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_10
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_559), .regcea(vdd), .wea(write_enable_22), .addra(address_22), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_13), .regceb(vdd), .web(write_enable_13), .addrb(address_13), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_566[131:131]), .sbiterrb(_566[130:130]), .doutb(_566[129:66]), .dbiterra(_566[65:65]), .sbiterra(_566[64:64]), .douta(_566[63:0]) );
    assign _567 = _566[63:0];
    assign _497 = ~ PHASE_4;
    assign _15 = _497;
    always @(posedge _84) begin
        if (_82)
            PHASE_4 <= _495;
        else
            if (_72)
                PHASE_4 <= _15;
    end
    assign _579 = PHASE_4 ? _578 : _567;
    assign address_23 = _764 ? _199 : _759;
    assign write_enable_23 = _757 & _764;
    assign address_24 = _764 ? _164 : _68;
    assign _766 = ~ _764;
    assign read_enable_19 = _752 & _766;
    assign _764 = ~ PHASE_7;
    assign write_enable_24 = _750 & _764;
    assign _768 = write_enable_24 | read_enable_19;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_11
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_768), .regcea(vdd), .wea(write_enable_24), .addra(address_24), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_23), .regceb(vdd), .web(write_enable_23), .addrb(address_23), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_773[131:131]), .sbiterrb(_773[130:130]), .doutb(_773[129:66]), .dbiterra(_773[65:65]), .sbiterra(_773[64:64]), .douta(_773[63:0]) );
    assign _774 = _773[63:0];
    assign address_25 = PHASE_7 ? _199 : _759;
    assign _757 = _129 & _720;
    assign write_enable_25 = _757 & PHASE_7;
    assign _682 = _674[129:66];
    assign _681 = _661[129:66];
    assign _683 = PHASE_5 ? _682 : _681;
    assign _679 = _619[129:66];
    assign _678 = _605[129:66];
    assign q1_1 = PHASE_6 ? _679 : _678;
    assign _684 = _586 ? _683 : q1_1;
    assign address_26 = _663 ? _657 : _656;
    assign _669 = ~ _663;
    assign read_enable_20 = _102 & _669;
    assign address_27 = _663 ? _60 : _639;
    assign _665 = ~ _663;
    assign read_enable_21 = _102 & _665;
    assign _663 = ~ PHASE_5;
    assign write_enable_27 = _622 & _663;
    assign _667 = write_enable_27 | read_enable_21;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_12
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_667), .regcea(vdd), .wea(write_enable_27), .addra(address_27), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_20), .regceb(vdd), .web(write_enable_26), .addrb(address_26), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_674[131:131]), .sbiterrb(_674[130:130]), .doutb(_674[129:66]), .dbiterra(_674[65:65]), .sbiterra(_674[64:64]), .douta(_674[63:0]) );
    assign _675 = _674[63:0];
    assign _655 = _172[11:11];
    assign _654 = _172[10:10];
    assign _653 = _172[9:9];
    assign _652 = _172[8:8];
    assign _651 = _172[7:7];
    assign _650 = _172[6:6];
    assign _649 = _172[5:5];
    assign _648 = _172[4:4];
    assign _647 = _172[3:3];
    assign _646 = _172[2:2];
    assign _645 = _172[1:1];
    assign _644 = _172[0:0];
    assign _656 = { _644, _645, _646, _647, _648, _649, _650, _651, _652, _653, _654, _655 };
    assign address_28 = PHASE_5 ? _657 : _656;
    assign _641 = ~ PHASE_5;
    assign read_enable_22 = _102 & _641;
    assign data_25 = wr_d5;
    assign _638 = _137[11:11];
    assign _637 = _137[10:10];
    assign _636 = _137[9:9];
    assign _635 = _137[8:8];
    assign _634 = _137[7:7];
    assign _633 = _137[6:6];
    assign _632 = _137[5:5];
    assign _631 = _137[4:4];
    assign _630 = _137[3:3];
    assign _629 = _137[2:2];
    assign _628 = _137[1:1];
    assign _627 = _137[0:0];
    assign _639 = { _627, _628, _629, _630, _631, _632, _633, _634, _635, _636, _637, _638 };
    assign address_29 = PHASE_5 ? _60 : _639;
    assign _624 = ~ PHASE_5;
    assign read_enable_23 = _102 & _624;
    assign _622 = _62[5:5];
    assign write_enable_29 = _622 & PHASE_5;
    assign _626 = write_enable_29 | read_enable_23;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_13
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_626), .regcea(vdd), .wea(write_enable_29), .addra(address_29), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_22), .regceb(vdd), .web(write_enable_28), .addrb(address_28), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_661[131:131]), .sbiterrb(_661[130:130]), .doutb(_661[129:66]), .dbiterra(_661[65:65]), .sbiterra(_661[64:64]), .douta(_661[63:0]) );
    assign _662 = _661[63:0];
    assign _583 = ~ PHASE_5;
    assign _19 = _583;
    always @(posedge _84) begin
        if (_82)
            PHASE_5 <= _581;
        else
            if (_72)
                PHASE_5 <= _19;
    end
    assign _676 = PHASE_5 ? _675 : _662;
    assign address_30 = _607 ? _199 : _172;
    assign _614 = ~ _607;
    assign read_enable_24 = _102 & _614;
    assign write_enable_30 = _598 & _607;
    assign _616 = write_enable_30 | read_enable_24;
    assign address_31 = _607 ? _164 : _137;
    assign _609 = ~ _607;
    assign read_enable_25 = _102 & _609;
    assign _607 = ~ PHASE_6;
    assign write_enable_31 = _591 & _607;
    assign _611 = write_enable_31 | read_enable_25;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_14
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_611), .regcea(vdd), .wea(write_enable_31), .addra(address_31), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_616), .regceb(vdd), .web(write_enable_30), .addrb(address_30), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_619[131:131]), .sbiterrb(_619[130:130]), .doutb(_619[129:66]), .dbiterra(_619[65:65]), .sbiterra(_619[64:64]), .douta(_619[63:0]) );
    assign _620 = _619[63:0];
    assign _687 = _686[127:64];
    assign data_27 = _687;
    assign address_32 = PHASE_6 ? _199 : _172;
    assign _600 = ~ PHASE_6;
    assign read_enable_26 = _102 & _600;
    assign _597 = ~ _130;
    assign _598 = _129 & _597;
    assign write_enable_32 = _598 & PHASE_6;
    assign _602 = write_enable_32 | read_enable_26;
    assign address_33 = PHASE_6 ? _164 : _137;
    assign _593 = ~ PHASE_6;
    assign read_enable_27 = _102 & _593;
    assign _590 = ~ _130;
    assign _591 = _129 & _590;
    assign write_enable_33 = _591 & PHASE_6;
    assign _595 = write_enable_33 | read_enable_27;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_15
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_595), .regcea(vdd), .wea(write_enable_33), .addra(address_33), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_602), .regceb(vdd), .web(write_enable_32), .addrb(address_32), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_605[131:131]), .sbiterrb(_605[130:130]), .doutb(_605[129:66]), .dbiterra(_605[65:65]), .sbiterra(_605[64:64]), .douta(_605[63:0]) );
    assign _606 = _605[63:0];
    assign _688 = ~ PHASE_6;
    assign _21 = _688;
    always @(posedge _84) begin
        if (_82)
            PHASE_6 <= _588;
        else
            if (_99)
                PHASE_6 <= _21;
    end
    assign q0_1 = PHASE_6 ? _620 : _606;
    always @(posedge _84) begin
        if (_82)
            _586 <= _585;
        else
            _586 <= _92;
    end
    assign _677 = _586 ? _676 : q0_1;
    dp_36
        dp_4
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_677), .d2(_684), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_686[191:128]), .q2(_686[127:64]), .q1(_686[63:0]) );
    assign _689 = _686[63:0];
    assign data_31 = _689;
    assign address_34 = PHASE_7 ? _164 : _68;
    assign _753 = ~ PHASE_7;
    assign _752 = _70[5:5];
    assign read_enable_28 = _752 & _753;
    always @(posedge _84) begin
        if (_82)
            _723 <= _722;
        else
            _723 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _726 <= _725;
        else
            _726 <= _723;
    end
    always @(posedge _84) begin
        if (_82)
            _729 <= _728;
        else
            _729 <= _726;
    end
    always @(posedge _84) begin
        if (_82)
            _732 <= _731;
        else
            _732 <= _729;
    end
    always @(posedge _84) begin
        if (_82)
            _735 <= _734;
        else
            _735 <= _732;
    end
    always @(posedge _84) begin
        if (_82)
            _738 <= _737;
        else
            _738 <= _735;
    end
    always @(posedge _84) begin
        if (_82)
            _741 <= _740;
        else
            _741 <= _738;
    end
    always @(posedge _84) begin
        if (_82)
            _744 <= _743;
        else
            _744 <= _741;
    end
    always @(posedge _84) begin
        if (_82)
            _747 <= _746;
        else
            _747 <= _744;
    end
    assign _748 = ~ _747;
    always @(posedge _84) begin
        if (_82)
            _696 <= _695;
        else
            _696 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _699 <= _698;
        else
            _699 <= _696;
    end
    always @(posedge _84) begin
        if (_82)
            _702 <= _701;
        else
            _702 <= _699;
    end
    always @(posedge _84) begin
        if (_82)
            _705 <= _704;
        else
            _705 <= _702;
    end
    always @(posedge _84) begin
        if (_82)
            _708 <= _707;
        else
            _708 <= _705;
    end
    always @(posedge _84) begin
        if (_82)
            _711 <= _710;
        else
            _711 <= _708;
    end
    always @(posedge _84) begin
        if (_82)
            _714 <= _713;
        else
            _714 <= _711;
    end
    always @(posedge _84) begin
        if (_82)
            _717 <= _716;
        else
            _717 <= _714;
    end
    always @(posedge _84) begin
        if (_82)
            _720 <= _719;
        else
            _720 <= _717;
    end
    assign _749 = _720 & _748;
    assign _750 = _129 & _749;
    assign write_enable_34 = _750 & PHASE_7;
    assign _755 = write_enable_34 | read_enable_28;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_16
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_755), .regcea(vdd), .wea(write_enable_34), .addra(address_34), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_25), .regceb(vdd), .web(write_enable_25), .addrb(address_25), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_762[131:131]), .sbiterrb(_762[130:130]), .doutb(_762[129:66]), .dbiterra(_762[65:65]), .sbiterra(_762[64:64]), .douta(_762[63:0]) );
    assign _763 = _762[63:0];
    assign _693 = ~ PHASE_7;
    assign _23 = _693;
    always @(posedge _84) begin
        if (_82)
            PHASE_7 <= _691;
        else
            if (_72)
                PHASE_7 <= _23;
    end
    assign _775 = PHASE_7 ? _774 : _763;
    assign address_35 = _960 ? _199 : _955;
    assign write_enable_35 = _953 & _960;
    assign address_36 = _960 ? _164 : _68;
    assign _962 = ~ _960;
    assign read_enable_29 = _948 & _962;
    assign _960 = ~ PHASE_10;
    assign write_enable_36 = _946 & _960;
    assign _964 = write_enable_36 | read_enable_29;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_17
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_964), .regcea(vdd), .wea(write_enable_36), .addra(address_36), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_35), .regceb(vdd), .web(write_enable_35), .addrb(address_35), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_969[131:131]), .sbiterrb(_969[130:130]), .doutb(_969[129:66]), .dbiterra(_969[65:65]), .sbiterra(_969[64:64]), .douta(_969[63:0]) );
    assign _970 = _969[63:0];
    assign address_37 = PHASE_10 ? _199 : _955;
    assign _953 = _129 & _916;
    assign write_enable_37 = _953 & PHASE_10;
    assign _878 = _870[129:66];
    assign _877 = _857[129:66];
    assign _879 = PHASE_8 ? _878 : _877;
    assign _875 = _815[129:66];
    assign _874 = _801[129:66];
    assign q1_2 = PHASE_9 ? _875 : _874;
    assign _880 = _782 ? _879 : q1_2;
    assign address_38 = _859 ? _853 : _852;
    assign _865 = ~ _859;
    assign read_enable_30 = _102 & _865;
    assign address_39 = _859 ? _60 : _835;
    assign _861 = ~ _859;
    assign read_enable_31 = _102 & _861;
    assign _859 = ~ PHASE_8;
    assign write_enable_39 = _818 & _859;
    assign _863 = write_enable_39 | read_enable_31;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_18
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_863), .regcea(vdd), .wea(write_enable_39), .addra(address_39), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_30), .regceb(vdd), .web(write_enable_38), .addrb(address_38), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_870[131:131]), .sbiterrb(_870[130:130]), .doutb(_870[129:66]), .dbiterra(_870[65:65]), .sbiterra(_870[64:64]), .douta(_870[63:0]) );
    assign _871 = _870[63:0];
    assign _851 = _172[11:11];
    assign _850 = _172[10:10];
    assign _849 = _172[9:9];
    assign _848 = _172[8:8];
    assign _847 = _172[7:7];
    assign _846 = _172[6:6];
    assign _845 = _172[5:5];
    assign _844 = _172[4:4];
    assign _843 = _172[3:3];
    assign _842 = _172[2:2];
    assign _841 = _172[1:1];
    assign _840 = _172[0:0];
    assign _852 = { _840, _841, _842, _843, _844, _845, _846, _847, _848, _849, _850, _851 };
    assign address_40 = PHASE_8 ? _853 : _852;
    assign _837 = ~ PHASE_8;
    assign read_enable_32 = _102 & _837;
    assign data_37 = wr_d4;
    assign _834 = _137[11:11];
    assign _833 = _137[10:10];
    assign _832 = _137[9:9];
    assign _831 = _137[8:8];
    assign _830 = _137[7:7];
    assign _829 = _137[6:6];
    assign _828 = _137[5:5];
    assign _827 = _137[4:4];
    assign _826 = _137[3:3];
    assign _825 = _137[2:2];
    assign _824 = _137[1:1];
    assign _823 = _137[0:0];
    assign _835 = { _823, _824, _825, _826, _827, _828, _829, _830, _831, _832, _833, _834 };
    assign address_41 = PHASE_8 ? _60 : _835;
    assign _820 = ~ PHASE_8;
    assign read_enable_33 = _102 & _820;
    assign _818 = _62[4:4];
    assign write_enable_41 = _818 & PHASE_8;
    assign _822 = write_enable_41 | read_enable_33;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_19
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_822), .regcea(vdd), .wea(write_enable_41), .addra(address_41), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_32), .regceb(vdd), .web(write_enable_40), .addrb(address_40), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_857[131:131]), .sbiterrb(_857[130:130]), .doutb(_857[129:66]), .dbiterra(_857[65:65]), .sbiterra(_857[64:64]), .douta(_857[63:0]) );
    assign _858 = _857[63:0];
    assign _779 = ~ PHASE_8;
    assign _27 = _779;
    always @(posedge _84) begin
        if (_82)
            PHASE_8 <= _777;
        else
            if (_72)
                PHASE_8 <= _27;
    end
    assign _872 = PHASE_8 ? _871 : _858;
    assign address_42 = _803 ? _199 : _172;
    assign _810 = ~ _803;
    assign read_enable_34 = _102 & _810;
    assign write_enable_42 = _794 & _803;
    assign _812 = write_enable_42 | read_enable_34;
    assign address_43 = _803 ? _164 : _137;
    assign _805 = ~ _803;
    assign read_enable_35 = _102 & _805;
    assign _803 = ~ PHASE_9;
    assign write_enable_43 = _787 & _803;
    assign _807 = write_enable_43 | read_enable_35;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_20
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_807), .regcea(vdd), .wea(write_enable_43), .addra(address_43), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_812), .regceb(vdd), .web(write_enable_42), .addrb(address_42), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_815[131:131]), .sbiterrb(_815[130:130]), .doutb(_815[129:66]), .dbiterra(_815[65:65]), .sbiterra(_815[64:64]), .douta(_815[63:0]) );
    assign _816 = _815[63:0];
    assign _883 = _882[127:64];
    assign data_39 = _883;
    assign address_44 = PHASE_9 ? _199 : _172;
    assign _796 = ~ PHASE_9;
    assign read_enable_36 = _102 & _796;
    assign _793 = ~ _130;
    assign _794 = _129 & _793;
    assign write_enable_44 = _794 & PHASE_9;
    assign _798 = write_enable_44 | read_enable_36;
    assign address_45 = PHASE_9 ? _164 : _137;
    assign _789 = ~ PHASE_9;
    assign read_enable_37 = _102 & _789;
    assign _786 = ~ _130;
    assign _787 = _129 & _786;
    assign write_enable_45 = _787 & PHASE_9;
    assign _791 = write_enable_45 | read_enable_37;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_21
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_791), .regcea(vdd), .wea(write_enable_45), .addra(address_45), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_798), .regceb(vdd), .web(write_enable_44), .addrb(address_44), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_801[131:131]), .sbiterrb(_801[130:130]), .doutb(_801[129:66]), .dbiterra(_801[65:65]), .sbiterra(_801[64:64]), .douta(_801[63:0]) );
    assign _802 = _801[63:0];
    assign _884 = ~ PHASE_9;
    assign _29 = _884;
    always @(posedge _84) begin
        if (_82)
            PHASE_9 <= _784;
        else
            if (_99)
                PHASE_9 <= _29;
    end
    assign q0_2 = PHASE_9 ? _816 : _802;
    always @(posedge _84) begin
        if (_82)
            _782 <= _781;
        else
            _782 <= _92;
    end
    assign _873 = _782 ? _872 : q0_2;
    dp_35
        dp_3
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_873), .d2(_880), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_882[191:128]), .q2(_882[127:64]), .q1(_882[63:0]) );
    assign _885 = _882[63:0];
    assign data_43 = _885;
    assign address_46 = PHASE_10 ? _164 : _68;
    assign _949 = ~ PHASE_10;
    assign _948 = _70[4:4];
    assign read_enable_38 = _948 & _949;
    always @(posedge _84) begin
        if (_82)
            _919 <= _918;
        else
            _919 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _922 <= _921;
        else
            _922 <= _919;
    end
    always @(posedge _84) begin
        if (_82)
            _925 <= _924;
        else
            _925 <= _922;
    end
    always @(posedge _84) begin
        if (_82)
            _928 <= _927;
        else
            _928 <= _925;
    end
    always @(posedge _84) begin
        if (_82)
            _931 <= _930;
        else
            _931 <= _928;
    end
    always @(posedge _84) begin
        if (_82)
            _934 <= _933;
        else
            _934 <= _931;
    end
    always @(posedge _84) begin
        if (_82)
            _937 <= _936;
        else
            _937 <= _934;
    end
    always @(posedge _84) begin
        if (_82)
            _940 <= _939;
        else
            _940 <= _937;
    end
    always @(posedge _84) begin
        if (_82)
            _943 <= _942;
        else
            _943 <= _940;
    end
    assign _944 = ~ _943;
    always @(posedge _84) begin
        if (_82)
            _892 <= _891;
        else
            _892 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _895 <= _894;
        else
            _895 <= _892;
    end
    always @(posedge _84) begin
        if (_82)
            _898 <= _897;
        else
            _898 <= _895;
    end
    always @(posedge _84) begin
        if (_82)
            _901 <= _900;
        else
            _901 <= _898;
    end
    always @(posedge _84) begin
        if (_82)
            _904 <= _903;
        else
            _904 <= _901;
    end
    always @(posedge _84) begin
        if (_82)
            _907 <= _906;
        else
            _907 <= _904;
    end
    always @(posedge _84) begin
        if (_82)
            _910 <= _909;
        else
            _910 <= _907;
    end
    always @(posedge _84) begin
        if (_82)
            _913 <= _912;
        else
            _913 <= _910;
    end
    always @(posedge _84) begin
        if (_82)
            _916 <= _915;
        else
            _916 <= _913;
    end
    assign _945 = _916 & _944;
    assign _946 = _129 & _945;
    assign write_enable_46 = _946 & PHASE_10;
    assign _951 = write_enable_46 | read_enable_38;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_22
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_951), .regcea(vdd), .wea(write_enable_46), .addra(address_46), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_37), .regceb(vdd), .web(write_enable_37), .addrb(address_37), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_958[131:131]), .sbiterrb(_958[130:130]), .doutb(_958[129:66]), .dbiterra(_958[65:65]), .sbiterra(_958[64:64]), .douta(_958[63:0]) );
    assign _959 = _958[63:0];
    assign _889 = ~ PHASE_10;
    assign _31 = _889;
    always @(posedge _84) begin
        if (_82)
            PHASE_10 <= _887;
        else
            if (_72)
                PHASE_10 <= _31;
    end
    assign _971 = PHASE_10 ? _970 : _959;
    assign address_47 = _1156 ? _199 : _1151;
    assign write_enable_47 = _1149 & _1156;
    assign address_48 = _1156 ? _164 : _68;
    assign _1158 = ~ _1156;
    assign read_enable_39 = _1144 & _1158;
    assign _1156 = ~ PHASE_13;
    assign write_enable_48 = _1142 & _1156;
    assign _1160 = write_enable_48 | read_enable_39;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_23
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1160), .regcea(vdd), .wea(write_enable_48), .addra(address_48), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_47), .regceb(vdd), .web(write_enable_47), .addrb(address_47), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1165[131:131]), .sbiterrb(_1165[130:130]), .doutb(_1165[129:66]), .dbiterra(_1165[65:65]), .sbiterra(_1165[64:64]), .douta(_1165[63:0]) );
    assign _1166 = _1165[63:0];
    assign address_49 = PHASE_13 ? _199 : _1151;
    assign _1149 = _129 & _1112;
    assign write_enable_49 = _1149 & PHASE_13;
    assign _1074 = _1066[129:66];
    assign _1073 = _1053[129:66];
    assign _1075 = PHASE_11 ? _1074 : _1073;
    assign _1071 = _1011[129:66];
    assign _1070 = _997[129:66];
    assign q1_3 = PHASE_12 ? _1071 : _1070;
    assign _1076 = _978 ? _1075 : q1_3;
    assign address_50 = _1055 ? _1049 : _1048;
    assign _1061 = ~ _1055;
    assign read_enable_40 = _102 & _1061;
    assign address_51 = _1055 ? _60 : _1031;
    assign _1057 = ~ _1055;
    assign read_enable_41 = _102 & _1057;
    assign _1055 = ~ PHASE_11;
    assign write_enable_51 = _1014 & _1055;
    assign _1059 = write_enable_51 | read_enable_41;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_24
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1059), .regcea(vdd), .wea(write_enable_51), .addra(address_51), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_40), .regceb(vdd), .web(write_enable_50), .addrb(address_50), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1066[131:131]), .sbiterrb(_1066[130:130]), .doutb(_1066[129:66]), .dbiterra(_1066[65:65]), .sbiterra(_1066[64:64]), .douta(_1066[63:0]) );
    assign _1067 = _1066[63:0];
    assign _1047 = _172[11:11];
    assign _1046 = _172[10:10];
    assign _1045 = _172[9:9];
    assign _1044 = _172[8:8];
    assign _1043 = _172[7:7];
    assign _1042 = _172[6:6];
    assign _1041 = _172[5:5];
    assign _1040 = _172[4:4];
    assign _1039 = _172[3:3];
    assign _1038 = _172[2:2];
    assign _1037 = _172[1:1];
    assign _1036 = _172[0:0];
    assign _1048 = { _1036, _1037, _1038, _1039, _1040, _1041, _1042, _1043, _1044, _1045, _1046, _1047 };
    assign address_52 = PHASE_11 ? _1049 : _1048;
    assign _1033 = ~ PHASE_11;
    assign read_enable_42 = _102 & _1033;
    assign data_49 = wr_d3;
    assign _1030 = _137[11:11];
    assign _1029 = _137[10:10];
    assign _1028 = _137[9:9];
    assign _1027 = _137[8:8];
    assign _1026 = _137[7:7];
    assign _1025 = _137[6:6];
    assign _1024 = _137[5:5];
    assign _1023 = _137[4:4];
    assign _1022 = _137[3:3];
    assign _1021 = _137[2:2];
    assign _1020 = _137[1:1];
    assign _1019 = _137[0:0];
    assign _1031 = { _1019, _1020, _1021, _1022, _1023, _1024, _1025, _1026, _1027, _1028, _1029, _1030 };
    assign address_53 = PHASE_11 ? _60 : _1031;
    assign _1016 = ~ PHASE_11;
    assign read_enable_43 = _102 & _1016;
    assign _1014 = _62[3:3];
    assign write_enable_53 = _1014 & PHASE_11;
    assign _1018 = write_enable_53 | read_enable_43;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_25
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1018), .regcea(vdd), .wea(write_enable_53), .addra(address_53), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_42), .regceb(vdd), .web(write_enable_52), .addrb(address_52), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1053[131:131]), .sbiterrb(_1053[130:130]), .doutb(_1053[129:66]), .dbiterra(_1053[65:65]), .sbiterra(_1053[64:64]), .douta(_1053[63:0]) );
    assign _1054 = _1053[63:0];
    assign _975 = ~ PHASE_11;
    assign _35 = _975;
    always @(posedge _84) begin
        if (_82)
            PHASE_11 <= _973;
        else
            if (_72)
                PHASE_11 <= _35;
    end
    assign _1068 = PHASE_11 ? _1067 : _1054;
    assign address_54 = _999 ? _199 : _172;
    assign _1006 = ~ _999;
    assign read_enable_44 = _102 & _1006;
    assign write_enable_54 = _990 & _999;
    assign _1008 = write_enable_54 | read_enable_44;
    assign address_55 = _999 ? _164 : _137;
    assign _1001 = ~ _999;
    assign read_enable_45 = _102 & _1001;
    assign _999 = ~ PHASE_12;
    assign write_enable_55 = _983 & _999;
    assign _1003 = write_enable_55 | read_enable_45;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_26
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1003), .regcea(vdd), .wea(write_enable_55), .addra(address_55), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1008), .regceb(vdd), .web(write_enable_54), .addrb(address_54), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1011[131:131]), .sbiterrb(_1011[130:130]), .doutb(_1011[129:66]), .dbiterra(_1011[65:65]), .sbiterra(_1011[64:64]), .douta(_1011[63:0]) );
    assign _1012 = _1011[63:0];
    assign _1079 = _1078[127:64];
    assign data_51 = _1079;
    assign address_56 = PHASE_12 ? _199 : _172;
    assign _992 = ~ PHASE_12;
    assign read_enable_46 = _102 & _992;
    assign _989 = ~ _130;
    assign _990 = _129 & _989;
    assign write_enable_56 = _990 & PHASE_12;
    assign _994 = write_enable_56 | read_enable_46;
    assign address_57 = PHASE_12 ? _164 : _137;
    assign _985 = ~ PHASE_12;
    assign read_enable_47 = _102 & _985;
    assign _982 = ~ _130;
    assign _983 = _129 & _982;
    assign write_enable_57 = _983 & PHASE_12;
    assign _987 = write_enable_57 | read_enable_47;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_27
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_987), .regcea(vdd), .wea(write_enable_57), .addra(address_57), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_994), .regceb(vdd), .web(write_enable_56), .addrb(address_56), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_997[131:131]), .sbiterrb(_997[130:130]), .doutb(_997[129:66]), .dbiterra(_997[65:65]), .sbiterra(_997[64:64]), .douta(_997[63:0]) );
    assign _998 = _997[63:0];
    assign _1080 = ~ PHASE_12;
    assign _37 = _1080;
    always @(posedge _84) begin
        if (_82)
            PHASE_12 <= _980;
        else
            if (_99)
                PHASE_12 <= _37;
    end
    assign q0_3 = PHASE_12 ? _1012 : _998;
    always @(posedge _84) begin
        if (_82)
            _978 <= _977;
        else
            _978 <= _92;
    end
    assign _1069 = _978 ? _1068 : q0_3;
    dp_34
        dp_2
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1069), .d2(_1076), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1078[191:128]), .q2(_1078[127:64]), .q1(_1078[63:0]) );
    assign _1081 = _1078[63:0];
    assign data_55 = _1081;
    assign address_58 = PHASE_13 ? _164 : _68;
    assign _1145 = ~ PHASE_13;
    assign _1144 = _70[3:3];
    assign read_enable_48 = _1144 & _1145;
    always @(posedge _84) begin
        if (_82)
            _1115 <= _1114;
        else
            _1115 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1118 <= _1117;
        else
            _1118 <= _1115;
    end
    always @(posedge _84) begin
        if (_82)
            _1121 <= _1120;
        else
            _1121 <= _1118;
    end
    always @(posedge _84) begin
        if (_82)
            _1124 <= _1123;
        else
            _1124 <= _1121;
    end
    always @(posedge _84) begin
        if (_82)
            _1127 <= _1126;
        else
            _1127 <= _1124;
    end
    always @(posedge _84) begin
        if (_82)
            _1130 <= _1129;
        else
            _1130 <= _1127;
    end
    always @(posedge _84) begin
        if (_82)
            _1133 <= _1132;
        else
            _1133 <= _1130;
    end
    always @(posedge _84) begin
        if (_82)
            _1136 <= _1135;
        else
            _1136 <= _1133;
    end
    always @(posedge _84) begin
        if (_82)
            _1139 <= _1138;
        else
            _1139 <= _1136;
    end
    assign _1140 = ~ _1139;
    always @(posedge _84) begin
        if (_82)
            _1088 <= _1087;
        else
            _1088 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1091 <= _1090;
        else
            _1091 <= _1088;
    end
    always @(posedge _84) begin
        if (_82)
            _1094 <= _1093;
        else
            _1094 <= _1091;
    end
    always @(posedge _84) begin
        if (_82)
            _1097 <= _1096;
        else
            _1097 <= _1094;
    end
    always @(posedge _84) begin
        if (_82)
            _1100 <= _1099;
        else
            _1100 <= _1097;
    end
    always @(posedge _84) begin
        if (_82)
            _1103 <= _1102;
        else
            _1103 <= _1100;
    end
    always @(posedge _84) begin
        if (_82)
            _1106 <= _1105;
        else
            _1106 <= _1103;
    end
    always @(posedge _84) begin
        if (_82)
            _1109 <= _1108;
        else
            _1109 <= _1106;
    end
    always @(posedge _84) begin
        if (_82)
            _1112 <= _1111;
        else
            _1112 <= _1109;
    end
    assign _1141 = _1112 & _1140;
    assign _1142 = _129 & _1141;
    assign write_enable_58 = _1142 & PHASE_13;
    assign _1147 = write_enable_58 | read_enable_48;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_28
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1147), .regcea(vdd), .wea(write_enable_58), .addra(address_58), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_49), .regceb(vdd), .web(write_enable_49), .addrb(address_49), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1154[131:131]), .sbiterrb(_1154[130:130]), .doutb(_1154[129:66]), .dbiterra(_1154[65:65]), .sbiterra(_1154[64:64]), .douta(_1154[63:0]) );
    assign _1155 = _1154[63:0];
    assign _1085 = ~ PHASE_13;
    assign _39 = _1085;
    always @(posedge _84) begin
        if (_82)
            PHASE_13 <= _1083;
        else
            if (_72)
                PHASE_13 <= _39;
    end
    assign _1167 = PHASE_13 ? _1166 : _1155;
    assign address_59 = _1352 ? _199 : _1347;
    assign write_enable_59 = _1345 & _1352;
    assign address_60 = _1352 ? _164 : _68;
    assign _1354 = ~ _1352;
    assign read_enable_49 = _1340 & _1354;
    assign _1352 = ~ PHASE_16;
    assign write_enable_60 = _1338 & _1352;
    assign _1356 = write_enable_60 | read_enable_49;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_29
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1356), .regcea(vdd), .wea(write_enable_60), .addra(address_60), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_59), .regceb(vdd), .web(write_enable_59), .addrb(address_59), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1361[131:131]), .sbiterrb(_1361[130:130]), .doutb(_1361[129:66]), .dbiterra(_1361[65:65]), .sbiterra(_1361[64:64]), .douta(_1361[63:0]) );
    assign _1362 = _1361[63:0];
    assign address_61 = PHASE_16 ? _199 : _1347;
    assign _1345 = _129 & _1308;
    assign write_enable_61 = _1345 & PHASE_16;
    assign _1270 = _1262[129:66];
    assign _1269 = _1249[129:66];
    assign _1271 = PHASE_14 ? _1270 : _1269;
    assign _1267 = _1207[129:66];
    assign _1266 = _1193[129:66];
    assign q1_4 = PHASE_15 ? _1267 : _1266;
    assign _1272 = _1174 ? _1271 : q1_4;
    assign address_62 = _1251 ? _1245 : _1244;
    assign _1257 = ~ _1251;
    assign read_enable_50 = _102 & _1257;
    assign address_63 = _1251 ? _60 : _1227;
    assign _1253 = ~ _1251;
    assign read_enable_51 = _102 & _1253;
    assign _1251 = ~ PHASE_14;
    assign write_enable_63 = _1210 & _1251;
    assign _1255 = write_enable_63 | read_enable_51;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_30
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1255), .regcea(vdd), .wea(write_enable_63), .addra(address_63), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_50), .regceb(vdd), .web(write_enable_62), .addrb(address_62), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1262[131:131]), .sbiterrb(_1262[130:130]), .doutb(_1262[129:66]), .dbiterra(_1262[65:65]), .sbiterra(_1262[64:64]), .douta(_1262[63:0]) );
    assign _1263 = _1262[63:0];
    assign _1243 = _172[11:11];
    assign _1242 = _172[10:10];
    assign _1241 = _172[9:9];
    assign _1240 = _172[8:8];
    assign _1239 = _172[7:7];
    assign _1238 = _172[6:6];
    assign _1237 = _172[5:5];
    assign _1236 = _172[4:4];
    assign _1235 = _172[3:3];
    assign _1234 = _172[2:2];
    assign _1233 = _172[1:1];
    assign _1232 = _172[0:0];
    assign _1244 = { _1232, _1233, _1234, _1235, _1236, _1237, _1238, _1239, _1240, _1241, _1242, _1243 };
    assign address_64 = PHASE_14 ? _1245 : _1244;
    assign _1229 = ~ PHASE_14;
    assign read_enable_52 = _102 & _1229;
    assign data_61 = wr_d2;
    assign _1226 = _137[11:11];
    assign _1225 = _137[10:10];
    assign _1224 = _137[9:9];
    assign _1223 = _137[8:8];
    assign _1222 = _137[7:7];
    assign _1221 = _137[6:6];
    assign _1220 = _137[5:5];
    assign _1219 = _137[4:4];
    assign _1218 = _137[3:3];
    assign _1217 = _137[2:2];
    assign _1216 = _137[1:1];
    assign _1215 = _137[0:0];
    assign _1227 = { _1215, _1216, _1217, _1218, _1219, _1220, _1221, _1222, _1223, _1224, _1225, _1226 };
    assign address_65 = PHASE_14 ? _60 : _1227;
    assign _1212 = ~ PHASE_14;
    assign read_enable_53 = _102 & _1212;
    assign _1210 = _62[2:2];
    assign write_enable_65 = _1210 & PHASE_14;
    assign _1214 = write_enable_65 | read_enable_53;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_31
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1214), .regcea(vdd), .wea(write_enable_65), .addra(address_65), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_52), .regceb(vdd), .web(write_enable_64), .addrb(address_64), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1249[131:131]), .sbiterrb(_1249[130:130]), .doutb(_1249[129:66]), .dbiterra(_1249[65:65]), .sbiterra(_1249[64:64]), .douta(_1249[63:0]) );
    assign _1250 = _1249[63:0];
    assign _1171 = ~ PHASE_14;
    assign _43 = _1171;
    always @(posedge _84) begin
        if (_82)
            PHASE_14 <= _1169;
        else
            if (_72)
                PHASE_14 <= _43;
    end
    assign _1264 = PHASE_14 ? _1263 : _1250;
    assign address_66 = _1195 ? _199 : _172;
    assign _1202 = ~ _1195;
    assign read_enable_54 = _102 & _1202;
    assign write_enable_66 = _1186 & _1195;
    assign _1204 = write_enable_66 | read_enable_54;
    assign address_67 = _1195 ? _164 : _137;
    assign _1197 = ~ _1195;
    assign read_enable_55 = _102 & _1197;
    assign _1195 = ~ PHASE_15;
    assign write_enable_67 = _1179 & _1195;
    assign _1199 = write_enable_67 | read_enable_55;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_32
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1199), .regcea(vdd), .wea(write_enable_67), .addra(address_67), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1204), .regceb(vdd), .web(write_enable_66), .addrb(address_66), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1207[131:131]), .sbiterrb(_1207[130:130]), .doutb(_1207[129:66]), .dbiterra(_1207[65:65]), .sbiterra(_1207[64:64]), .douta(_1207[63:0]) );
    assign _1208 = _1207[63:0];
    assign _1275 = _1274[127:64];
    assign data_63 = _1275;
    assign address_68 = PHASE_15 ? _199 : _172;
    assign _1188 = ~ PHASE_15;
    assign read_enable_56 = _102 & _1188;
    assign _1185 = ~ _130;
    assign _1186 = _129 & _1185;
    assign write_enable_68 = _1186 & PHASE_15;
    assign _1190 = write_enable_68 | read_enable_56;
    assign address_69 = PHASE_15 ? _164 : _137;
    assign _1181 = ~ PHASE_15;
    assign read_enable_57 = _102 & _1181;
    assign _1178 = ~ _130;
    assign _1179 = _129 & _1178;
    assign write_enable_69 = _1179 & PHASE_15;
    assign _1183 = write_enable_69 | read_enable_57;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_33
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1183), .regcea(vdd), .wea(write_enable_69), .addra(address_69), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1190), .regceb(vdd), .web(write_enable_68), .addrb(address_68), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1193[131:131]), .sbiterrb(_1193[130:130]), .doutb(_1193[129:66]), .dbiterra(_1193[65:65]), .sbiterra(_1193[64:64]), .douta(_1193[63:0]) );
    assign _1194 = _1193[63:0];
    assign _1276 = ~ PHASE_15;
    assign _45 = _1276;
    always @(posedge _84) begin
        if (_82)
            PHASE_15 <= _1176;
        else
            if (_99)
                PHASE_15 <= _45;
    end
    assign q0_4 = PHASE_15 ? _1208 : _1194;
    always @(posedge _84) begin
        if (_82)
            _1174 <= _1173;
        else
            _1174 <= _92;
    end
    assign _1265 = _1174 ? _1264 : q0_4;
    dp_33
        dp_1
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1265), .d2(_1272), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1274[191:128]), .q2(_1274[127:64]), .q1(_1274[63:0]) );
    assign _1277 = _1274[63:0];
    assign data_67 = _1277;
    assign address_70 = PHASE_16 ? _164 : _68;
    assign _1341 = ~ PHASE_16;
    assign _1340 = _70[2:2];
    assign read_enable_58 = _1340 & _1341;
    always @(posedge _84) begin
        if (_82)
            _1311 <= _1310;
        else
            _1311 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1314 <= _1313;
        else
            _1314 <= _1311;
    end
    always @(posedge _84) begin
        if (_82)
            _1317 <= _1316;
        else
            _1317 <= _1314;
    end
    always @(posedge _84) begin
        if (_82)
            _1320 <= _1319;
        else
            _1320 <= _1317;
    end
    always @(posedge _84) begin
        if (_82)
            _1323 <= _1322;
        else
            _1323 <= _1320;
    end
    always @(posedge _84) begin
        if (_82)
            _1326 <= _1325;
        else
            _1326 <= _1323;
    end
    always @(posedge _84) begin
        if (_82)
            _1329 <= _1328;
        else
            _1329 <= _1326;
    end
    always @(posedge _84) begin
        if (_82)
            _1332 <= _1331;
        else
            _1332 <= _1329;
    end
    always @(posedge _84) begin
        if (_82)
            _1335 <= _1334;
        else
            _1335 <= _1332;
    end
    assign _1336 = ~ _1335;
    always @(posedge _84) begin
        if (_82)
            _1284 <= _1283;
        else
            _1284 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1287 <= _1286;
        else
            _1287 <= _1284;
    end
    always @(posedge _84) begin
        if (_82)
            _1290 <= _1289;
        else
            _1290 <= _1287;
    end
    always @(posedge _84) begin
        if (_82)
            _1293 <= _1292;
        else
            _1293 <= _1290;
    end
    always @(posedge _84) begin
        if (_82)
            _1296 <= _1295;
        else
            _1296 <= _1293;
    end
    always @(posedge _84) begin
        if (_82)
            _1299 <= _1298;
        else
            _1299 <= _1296;
    end
    always @(posedge _84) begin
        if (_82)
            _1302 <= _1301;
        else
            _1302 <= _1299;
    end
    always @(posedge _84) begin
        if (_82)
            _1305 <= _1304;
        else
            _1305 <= _1302;
    end
    always @(posedge _84) begin
        if (_82)
            _1308 <= _1307;
        else
            _1308 <= _1305;
    end
    assign _1337 = _1308 & _1336;
    assign _1338 = _129 & _1337;
    assign write_enable_70 = _1338 & PHASE_16;
    assign _1343 = write_enable_70 | read_enable_58;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_34
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1343), .regcea(vdd), .wea(write_enable_70), .addra(address_70), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_61), .regceb(vdd), .web(write_enable_61), .addrb(address_61), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1350[131:131]), .sbiterrb(_1350[130:130]), .doutb(_1350[129:66]), .dbiterra(_1350[65:65]), .sbiterra(_1350[64:64]), .douta(_1350[63:0]) );
    assign _1351 = _1350[63:0];
    assign _1281 = ~ PHASE_16;
    assign _47 = _1281;
    always @(posedge _84) begin
        if (_82)
            PHASE_16 <= _1279;
        else
            if (_72)
                PHASE_16 <= _47;
    end
    assign _1363 = PHASE_16 ? _1362 : _1351;
    assign address_71 = _1548 ? _199 : _1543;
    assign write_enable_71 = _1541 & _1548;
    assign address_72 = _1548 ? _164 : _68;
    assign _1550 = ~ _1548;
    assign read_enable_59 = _1536 & _1550;
    assign _1548 = ~ PHASE_19;
    assign write_enable_72 = _1534 & _1548;
    assign _1552 = write_enable_72 | read_enable_59;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_35
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1552), .regcea(vdd), .wea(write_enable_72), .addra(address_72), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_71), .regceb(vdd), .web(write_enable_71), .addrb(address_71), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1557[131:131]), .sbiterrb(_1557[130:130]), .doutb(_1557[129:66]), .dbiterra(_1557[65:65]), .sbiterra(_1557[64:64]), .douta(_1557[63:0]) );
    assign _1558 = _1557[63:0];
    assign address_73 = PHASE_19 ? _199 : _1543;
    assign _1541 = _129 & _1504;
    assign write_enable_73 = _1541 & PHASE_19;
    assign _1466 = _1458[129:66];
    assign _1465 = _1445[129:66];
    assign _1467 = PHASE_17 ? _1466 : _1465;
    assign _1463 = _1403[129:66];
    assign _1462 = _1389[129:66];
    assign q1_5 = PHASE_18 ? _1463 : _1462;
    assign _1468 = _1370 ? _1467 : q1_5;
    assign address_74 = _1447 ? _1441 : _1440;
    assign _1453 = ~ _1447;
    assign read_enable_60 = _102 & _1453;
    assign address_75 = _1447 ? _60 : _1423;
    assign _1449 = ~ _1447;
    assign read_enable_61 = _102 & _1449;
    assign _1447 = ~ PHASE_17;
    assign write_enable_75 = _1406 & _1447;
    assign _1451 = write_enable_75 | read_enable_61;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_36
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1451), .regcea(vdd), .wea(write_enable_75), .addra(address_75), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_60), .regceb(vdd), .web(write_enable_74), .addrb(address_74), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1458[131:131]), .sbiterrb(_1458[130:130]), .doutb(_1458[129:66]), .dbiterra(_1458[65:65]), .sbiterra(_1458[64:64]), .douta(_1458[63:0]) );
    assign _1459 = _1458[63:0];
    assign _1439 = _172[11:11];
    assign _1438 = _172[10:10];
    assign _1437 = _172[9:9];
    assign _1436 = _172[8:8];
    assign _1435 = _172[7:7];
    assign _1434 = _172[6:6];
    assign _1433 = _172[5:5];
    assign _1432 = _172[4:4];
    assign _1431 = _172[3:3];
    assign _1430 = _172[2:2];
    assign _1429 = _172[1:1];
    assign _1428 = _172[0:0];
    assign _1440 = { _1428, _1429, _1430, _1431, _1432, _1433, _1434, _1435, _1436, _1437, _1438, _1439 };
    assign address_76 = PHASE_17 ? _1441 : _1440;
    assign _1425 = ~ PHASE_17;
    assign read_enable_62 = _102 & _1425;
    assign data_73 = wr_d1;
    assign _1422 = _137[11:11];
    assign _1421 = _137[10:10];
    assign _1420 = _137[9:9];
    assign _1419 = _137[8:8];
    assign _1418 = _137[7:7];
    assign _1417 = _137[6:6];
    assign _1416 = _137[5:5];
    assign _1415 = _137[4:4];
    assign _1414 = _137[3:3];
    assign _1413 = _137[2:2];
    assign _1412 = _137[1:1];
    assign _1411 = _137[0:0];
    assign _1423 = { _1411, _1412, _1413, _1414, _1415, _1416, _1417, _1418, _1419, _1420, _1421, _1422 };
    assign address_77 = PHASE_17 ? _60 : _1423;
    assign _1408 = ~ PHASE_17;
    assign read_enable_63 = _102 & _1408;
    assign _1406 = _62[1:1];
    assign write_enable_77 = _1406 & PHASE_17;
    assign _1410 = write_enable_77 | read_enable_63;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_37
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1410), .regcea(vdd), .wea(write_enable_77), .addra(address_77), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_62), .regceb(vdd), .web(write_enable_76), .addrb(address_76), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1445[131:131]), .sbiterrb(_1445[130:130]), .doutb(_1445[129:66]), .dbiterra(_1445[65:65]), .sbiterra(_1445[64:64]), .douta(_1445[63:0]) );
    assign _1446 = _1445[63:0];
    assign _1367 = ~ PHASE_17;
    assign _51 = _1367;
    always @(posedge _84) begin
        if (_82)
            PHASE_17 <= _1365;
        else
            if (_72)
                PHASE_17 <= _51;
    end
    assign _1460 = PHASE_17 ? _1459 : _1446;
    assign address_78 = _1391 ? _199 : _172;
    assign _1398 = ~ _1391;
    assign read_enable_64 = _102 & _1398;
    assign write_enable_78 = _1382 & _1391;
    assign _1400 = write_enable_78 | read_enable_64;
    assign address_79 = _1391 ? _164 : _137;
    assign _1393 = ~ _1391;
    assign read_enable_65 = _102 & _1393;
    assign _1391 = ~ PHASE_18;
    assign write_enable_79 = _1375 & _1391;
    assign _1395 = write_enable_79 | read_enable_65;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_38
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1395), .regcea(vdd), .wea(write_enable_79), .addra(address_79), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1400), .regceb(vdd), .web(write_enable_78), .addrb(address_78), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1403[131:131]), .sbiterrb(_1403[130:130]), .doutb(_1403[129:66]), .dbiterra(_1403[65:65]), .sbiterra(_1403[64:64]), .douta(_1403[63:0]) );
    assign _1404 = _1403[63:0];
    assign _1471 = _1470[127:64];
    assign data_75 = _1471;
    assign address_80 = PHASE_18 ? _199 : _172;
    assign _1384 = ~ PHASE_18;
    assign read_enable_66 = _102 & _1384;
    assign _1381 = ~ _130;
    assign _1382 = _129 & _1381;
    assign write_enable_80 = _1382 & PHASE_18;
    assign _1386 = write_enable_80 | read_enable_66;
    assign address_81 = PHASE_18 ? _164 : _137;
    assign _1377 = ~ PHASE_18;
    assign read_enable_67 = _102 & _1377;
    assign _1374 = ~ _130;
    assign _1375 = _129 & _1374;
    assign write_enable_81 = _1375 & PHASE_18;
    assign _1379 = write_enable_81 | read_enable_67;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_39
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1379), .regcea(vdd), .wea(write_enable_81), .addra(address_81), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1386), .regceb(vdd), .web(write_enable_80), .addrb(address_80), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1389[131:131]), .sbiterrb(_1389[130:130]), .doutb(_1389[129:66]), .dbiterra(_1389[65:65]), .sbiterra(_1389[64:64]), .douta(_1389[63:0]) );
    assign _1390 = _1389[63:0];
    assign _1472 = ~ PHASE_18;
    assign _53 = _1472;
    always @(posedge _84) begin
        if (_82)
            PHASE_18 <= _1372;
        else
            if (_99)
                PHASE_18 <= _53;
    end
    assign q0_5 = PHASE_18 ? _1404 : _1390;
    always @(posedge _84) begin
        if (_82)
            _1370 <= _1369;
        else
            _1370 <= _92;
    end
    assign _1461 = _1370 ? _1460 : q0_5;
    dp_32
        dp_0
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1461), .d2(_1468), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1470[191:128]), .q2(_1470[127:64]), .q1(_1470[63:0]) );
    assign _1473 = _1470[63:0];
    assign data_79 = _1473;
    assign address_82 = PHASE_19 ? _164 : _68;
    assign _1537 = ~ PHASE_19;
    assign _1536 = _70[1:1];
    assign read_enable_68 = _1536 & _1537;
    always @(posedge _84) begin
        if (_82)
            _1507 <= _1506;
        else
            _1507 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1510 <= _1509;
        else
            _1510 <= _1507;
    end
    always @(posedge _84) begin
        if (_82)
            _1513 <= _1512;
        else
            _1513 <= _1510;
    end
    always @(posedge _84) begin
        if (_82)
            _1516 <= _1515;
        else
            _1516 <= _1513;
    end
    always @(posedge _84) begin
        if (_82)
            _1519 <= _1518;
        else
            _1519 <= _1516;
    end
    always @(posedge _84) begin
        if (_82)
            _1522 <= _1521;
        else
            _1522 <= _1519;
    end
    always @(posedge _84) begin
        if (_82)
            _1525 <= _1524;
        else
            _1525 <= _1522;
    end
    always @(posedge _84) begin
        if (_82)
            _1528 <= _1527;
        else
            _1528 <= _1525;
    end
    always @(posedge _84) begin
        if (_82)
            _1531 <= _1530;
        else
            _1531 <= _1528;
    end
    assign _1532 = ~ _1531;
    always @(posedge _84) begin
        if (_82)
            _1480 <= _1479;
        else
            _1480 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1483 <= _1482;
        else
            _1483 <= _1480;
    end
    always @(posedge _84) begin
        if (_82)
            _1486 <= _1485;
        else
            _1486 <= _1483;
    end
    always @(posedge _84) begin
        if (_82)
            _1489 <= _1488;
        else
            _1489 <= _1486;
    end
    always @(posedge _84) begin
        if (_82)
            _1492 <= _1491;
        else
            _1492 <= _1489;
    end
    always @(posedge _84) begin
        if (_82)
            _1495 <= _1494;
        else
            _1495 <= _1492;
    end
    always @(posedge _84) begin
        if (_82)
            _1498 <= _1497;
        else
            _1498 <= _1495;
    end
    always @(posedge _84) begin
        if (_82)
            _1501 <= _1500;
        else
            _1501 <= _1498;
    end
    always @(posedge _84) begin
        if (_82)
            _1504 <= _1503;
        else
            _1504 <= _1501;
    end
    assign _1533 = _1504 & _1532;
    assign _1534 = _129 & _1533;
    assign write_enable_82 = _1534 & PHASE_19;
    assign _1539 = write_enable_82 | read_enable_68;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_40
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1539), .regcea(vdd), .wea(write_enable_82), .addra(address_82), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_73), .regceb(vdd), .web(write_enable_73), .addrb(address_73), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1546[131:131]), .sbiterrb(_1546[130:130]), .doutb(_1546[129:66]), .dbiterra(_1546[65:65]), .sbiterra(_1546[64:64]), .douta(_1546[63:0]) );
    assign _1547 = _1546[63:0];
    assign _1477 = ~ PHASE_19;
    assign _55 = _1477;
    always @(posedge _84) begin
        if (_82)
            PHASE_19 <= _1475;
        else
            if (_72)
                PHASE_19 <= _55;
    end
    assign _1559 = PHASE_19 ? _1558 : _1547;
    assign address_83 = _1744 ? _199 : _1739;
    assign write_enable_83 = _1737 & _1744;
    assign address_84 = _1744 ? _164 : _68;
    assign _1746 = ~ _1744;
    assign read_enable_69 = _1732 & _1746;
    assign _1744 = ~ PHASE_22;
    assign write_enable_84 = _1730 & _1744;
    assign _1748 = write_enable_84 | read_enable_69;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_41
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1748), .regcea(vdd), .wea(write_enable_84), .addra(address_84), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_83), .regceb(vdd), .web(write_enable_83), .addrb(address_83), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1753[131:131]), .sbiterrb(_1753[130:130]), .doutb(_1753[129:66]), .dbiterra(_1753[65:65]), .sbiterra(_1753[64:64]), .douta(_1753[63:0]) );
    assign _1754 = _1753[63:0];
    assign address_85 = PHASE_22 ? _199 : _1739;
    assign _1737 = _129 & _1700;
    assign write_enable_85 = _1737 & PHASE_22;
    assign _292 = _91[521:518];
    assign _291 = _91[517:517];
    assign _289 = _91[513:513];
    assign _288 = _91[512:449];
    assign _287 = _91[448:385];
    assign _286 = _91[384:321];
    assign _285 = _91[320:257];
    assign _284 = _91[256:193];
    assign _283 = _91[192:129];
    assign _282 = _91[128:65];
    assign _1662 = _1654[129:66];
    assign _1661 = _1641[129:66];
    assign _1663 = PHASE_20 ? _1662 : _1661;
    assign _1659 = _1599[129:66];
    assign _1658 = _1585[129:66];
    assign q1_6 = PHASE_21 ? _1659 : _1658;
    assign _1664 = _1566 ? _1663 : q1_6;
    assign address_86 = _1643 ? _1637 : _1636;
    assign _1649 = ~ _1643;
    assign read_enable_70 = _102 & _1649;
    assign address_87 = _1643 ? _60 : _1619;
    assign _1645 = ~ _1643;
    assign read_enable_71 = _102 & _1645;
    assign _1643 = ~ PHASE_20;
    assign write_enable_87 = _1602 & _1643;
    assign _1647 = write_enable_87 | read_enable_71;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_42
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1647), .regcea(vdd), .wea(write_enable_87), .addra(address_87), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_70), .regceb(vdd), .web(write_enable_86), .addrb(address_86), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1654[131:131]), .sbiterrb(_1654[130:130]), .doutb(_1654[129:66]), .dbiterra(_1654[65:65]), .sbiterra(_1654[64:64]), .douta(_1654[63:0]) );
    assign _1655 = _1654[63:0];
    assign _1635 = _172[11:11];
    assign _1634 = _172[10:10];
    assign _1633 = _172[9:9];
    assign _1632 = _172[8:8];
    assign _1631 = _172[7:7];
    assign _1630 = _172[6:6];
    assign _1629 = _172[5:5];
    assign _1628 = _172[4:4];
    assign _1627 = _172[3:3];
    assign _1626 = _172[2:2];
    assign _1625 = _172[1:1];
    assign _1624 = _172[0:0];
    assign _1636 = { _1624, _1625, _1626, _1627, _1628, _1629, _1630, _1631, _1632, _1633, _1634, _1635 };
    assign address_88 = PHASE_20 ? _1637 : _1636;
    assign _1621 = ~ PHASE_20;
    assign read_enable_72 = _102 & _1621;
    assign data_85 = wr_d0;
    assign _60 = wr_addr;
    assign _1618 = _137[11:11];
    assign _1617 = _137[10:10];
    assign _1616 = _137[9:9];
    assign _1615 = _137[8:8];
    assign _1614 = _137[7:7];
    assign _1613 = _137[6:6];
    assign _1612 = _137[5:5];
    assign _1611 = _137[4:4];
    assign _1610 = _137[3:3];
    assign _1609 = _137[2:2];
    assign _1608 = _137[1:1];
    assign _1607 = _137[0:0];
    assign _1619 = { _1607, _1608, _1609, _1610, _1611, _1612, _1613, _1614, _1615, _1616, _1617, _1618 };
    assign address_89 = PHASE_20 ? _60 : _1619;
    assign _1604 = ~ PHASE_20;
    assign read_enable_73 = _102 & _1604;
    assign _62 = wr_en;
    assign _1602 = _62[0:0];
    assign write_enable_89 = _1602 & PHASE_20;
    assign _1606 = write_enable_89 | read_enable_73;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_43
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1606), .regcea(vdd), .wea(write_enable_89), .addra(address_89), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_72), .regceb(vdd), .web(write_enable_88), .addrb(address_88), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1641[131:131]), .sbiterrb(_1641[130:130]), .doutb(_1641[129:66]), .dbiterra(_1641[65:65]), .sbiterra(_1641[64:64]), .douta(_1641[63:0]) );
    assign _1642 = _1641[63:0];
    assign _1563 = ~ PHASE_20;
    assign _63 = _1563;
    always @(posedge _84) begin
        if (_82)
            PHASE_20 <= _1561;
        else
            if (_72)
                PHASE_20 <= _63;
    end
    assign _1656 = PHASE_20 ? _1655 : _1642;
    assign address_90 = _1587 ? _199 : _172;
    assign _1594 = ~ _1587;
    assign read_enable_74 = _102 & _1594;
    assign write_enable_90 = _1578 & _1587;
    assign _1596 = write_enable_90 | read_enable_74;
    assign address_91 = _1587 ? _164 : _137;
    assign _1589 = ~ _1587;
    assign read_enable_75 = _102 & _1589;
    assign _1587 = ~ PHASE_21;
    assign write_enable_91 = _1571 & _1587;
    assign _1591 = write_enable_91 | read_enable_75;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_44
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1591), .regcea(vdd), .wea(write_enable_91), .addra(address_91), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1596), .regceb(vdd), .web(write_enable_90), .addrb(address_90), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1599[131:131]), .sbiterrb(_1599[130:130]), .doutb(_1599[129:66]), .dbiterra(_1599[65:65]), .sbiterra(_1599[64:64]), .douta(_1599[63:0]) );
    assign _1600 = _1599[63:0];
    assign _1667 = _1666[127:64];
    assign data_87 = _1667;
    always @(posedge _84) begin
        if (_82)
            _175 <= _174;
        else
            _175 <= _172;
    end
    always @(posedge _84) begin
        if (_82)
            _178 <= _177;
        else
            _178 <= _175;
    end
    always @(posedge _84) begin
        if (_82)
            _181 <= _180;
        else
            _181 <= _178;
    end
    always @(posedge _84) begin
        if (_82)
            _184 <= _183;
        else
            _184 <= _181;
    end
    always @(posedge _84) begin
        if (_82)
            _187 <= _186;
        else
            _187 <= _184;
    end
    always @(posedge _84) begin
        if (_82)
            _190 <= _189;
        else
            _190 <= _187;
    end
    always @(posedge _84) begin
        if (_82)
            _193 <= _192;
        else
            _193 <= _190;
    end
    always @(posedge _84) begin
        if (_82)
            _196 <= _195;
        else
            _196 <= _193;
    end
    always @(posedge _84) begin
        if (_82)
            _199 <= _198;
        else
            _199 <= _196;
    end
    assign _172 = _91[64:53];
    assign address_92 = PHASE_21 ? _199 : _172;
    assign _1580 = ~ PHASE_21;
    assign read_enable_76 = _102 & _1580;
    assign _1577 = ~ _130;
    assign _1578 = _129 & _1577;
    assign write_enable_92 = _1578 & PHASE_21;
    assign _1582 = write_enable_92 | read_enable_76;
    assign address_93 = PHASE_21 ? _164 : _137;
    assign _1573 = ~ PHASE_21;
    assign read_enable_77 = _102 & _1573;
    assign _1570 = ~ _130;
    assign _1571 = _129 & _1570;
    assign write_enable_93 = _1571 & PHASE_21;
    assign _1575 = write_enable_93 | read_enable_77;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_45
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1575), .regcea(vdd), .wea(write_enable_93), .addra(address_93), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1582), .regceb(vdd), .web(write_enable_92), .addrb(address_92), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1585[131:131]), .sbiterrb(_1585[130:130]), .doutb(_1585[129:66]), .dbiterra(_1585[65:65]), .sbiterra(_1585[64:64]), .douta(_1585[63:0]) );
    assign _1586 = _1585[63:0];
    assign _99 = _91[523:523];
    assign _1668 = ~ PHASE_21;
    assign _65 = _1668;
    always @(posedge _84) begin
        if (_82)
            PHASE_21 <= _1568;
        else
            if (_99)
                PHASE_21 <= _65;
    end
    assign q0_6 = PHASE_21 ? _1600 : _1586;
    assign _92 = _91[514:514];
    always @(posedge _84) begin
        if (_82)
            _1566 <= _1565;
        else
            _1566 <= _92;
    end
    assign _1657 = _1566 ? _1656 : q0_6;
    dp_31
        dp
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1657), .d2(_1664), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1666[191:128]), .q2(_1666[127:64]), .q1(_1666[63:0]) );
    assign _1669 = _1666[63:0];
    assign data_91 = _1669;
    assign _137 = _91[52:41];
    always @(posedge _84) begin
        if (_82)
            _140 <= _139;
        else
            _140 <= _137;
    end
    always @(posedge _84) begin
        if (_82)
            _143 <= _142;
        else
            _143 <= _140;
    end
    always @(posedge _84) begin
        if (_82)
            _146 <= _145;
        else
            _146 <= _143;
    end
    always @(posedge _84) begin
        if (_82)
            _149 <= _148;
        else
            _149 <= _146;
    end
    always @(posedge _84) begin
        if (_82)
            _152 <= _151;
        else
            _152 <= _149;
    end
    always @(posedge _84) begin
        if (_82)
            _155 <= _154;
        else
            _155 <= _152;
    end
    always @(posedge _84) begin
        if (_82)
            _158 <= _157;
        else
            _158 <= _155;
    end
    always @(posedge _84) begin
        if (_82)
            _161 <= _160;
        else
            _161 <= _158;
    end
    always @(posedge _84) begin
        if (_82)
            _164 <= _163;
        else
            _164 <= _161;
    end
    assign _68 = rd_addr;
    assign address_94 = PHASE_22 ? _164 : _68;
    assign _1733 = ~ PHASE_22;
    assign _70 = rd_en;
    assign _1732 = _70[0:0];
    assign read_enable_78 = _1732 & _1733;
    assign _290 = _91[516:516];
    always @(posedge _84) begin
        if (_82)
            _1703 <= _1702;
        else
            _1703 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1706 <= _1705;
        else
            _1706 <= _1703;
    end
    always @(posedge _84) begin
        if (_82)
            _1709 <= _1708;
        else
            _1709 <= _1706;
    end
    always @(posedge _84) begin
        if (_82)
            _1712 <= _1711;
        else
            _1712 <= _1709;
    end
    always @(posedge _84) begin
        if (_82)
            _1715 <= _1714;
        else
            _1715 <= _1712;
    end
    always @(posedge _84) begin
        if (_82)
            _1718 <= _1717;
        else
            _1718 <= _1715;
    end
    always @(posedge _84) begin
        if (_82)
            _1721 <= _1720;
        else
            _1721 <= _1718;
    end
    always @(posedge _84) begin
        if (_82)
            _1724 <= _1723;
        else
            _1724 <= _1721;
    end
    always @(posedge _84) begin
        if (_82)
            _1727 <= _1726;
        else
            _1727 <= _1724;
    end
    assign _1728 = ~ _1727;
    assign _130 = _91[515:515];
    always @(posedge _84) begin
        if (_82)
            _1676 <= _1675;
        else
            _1676 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1679 <= _1678;
        else
            _1679 <= _1676;
    end
    always @(posedge _84) begin
        if (_82)
            _1682 <= _1681;
        else
            _1682 <= _1679;
    end
    always @(posedge _84) begin
        if (_82)
            _1685 <= _1684;
        else
            _1685 <= _1682;
    end
    always @(posedge _84) begin
        if (_82)
            _1688 <= _1687;
        else
            _1688 <= _1685;
    end
    always @(posedge _84) begin
        if (_82)
            _1691 <= _1690;
        else
            _1691 <= _1688;
    end
    always @(posedge _84) begin
        if (_82)
            _1694 <= _1693;
        else
            _1694 <= _1691;
    end
    always @(posedge _84) begin
        if (_82)
            _1697 <= _1696;
        else
            _1697 <= _1694;
    end
    always @(posedge _84) begin
        if (_82)
            _1700 <= _1699;
        else
            _1700 <= _1697;
    end
    assign _1729 = _1700 & _1728;
    assign _102 = _91[522:522];
    always @(posedge _84) begin
        if (_82)
            _105 <= _104;
        else
            _105 <= _102;
    end
    always @(posedge _84) begin
        if (_82)
            _108 <= _107;
        else
            _108 <= _105;
    end
    always @(posedge _84) begin
        if (_82)
            _111 <= _110;
        else
            _111 <= _108;
    end
    always @(posedge _84) begin
        if (_82)
            _114 <= _113;
        else
            _114 <= _111;
    end
    always @(posedge _84) begin
        if (_82)
            _117 <= _116;
        else
            _117 <= _114;
    end
    always @(posedge _84) begin
        if (_82)
            _120 <= _119;
        else
            _120 <= _117;
    end
    always @(posedge _84) begin
        if (_82)
            _123 <= _122;
        else
            _123 <= _120;
    end
    always @(posedge _84) begin
        if (_82)
            _126 <= _125;
        else
            _126 <= _123;
    end
    always @(posedge _84) begin
        if (_82)
            _129 <= _128;
        else
            _129 <= _126;
    end
    assign _1730 = _129 & _1729;
    assign write_enable_94 = _1730 & PHASE_22;
    assign _1735 = write_enable_94 | read_enable_78;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_46
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1735), .regcea(vdd), .wea(write_enable_94), .addra(address_94), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_85), .regceb(vdd), .web(write_enable_85), .addrb(address_85), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1742[131:131]), .sbiterrb(_1742[130:130]), .doutb(_1742[129:66]), .dbiterra(_1742[65:65]), .sbiterra(_1742[64:64]), .douta(_1742[63:0]) );
    assign _1743 = _1742[63:0];
    assign _72 = flip;
    assign _1673 = ~ PHASE_22;
    assign _73 = _1673;
    always @(posedge _84) begin
        if (_82)
            PHASE_22 <= _1671;
        else
            if (_72)
                PHASE_22 <= _73;
    end
    assign _1755 = PHASE_22 ? _1754 : _1743;
    assign _76 = first_4step_pass;
    assign _78 = first_iter;
    assign _80 = start;
    assign _82 = clear;
    assign _84 = clock;
    ctrl
        ctrl
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .first_4step_pass(_76), .flip(_91[523:523]), .read_write_enable(_91[522:522]), .index(_91[521:518]), .valid(_91[517:517]), .twiddle_stage(_91[516:516]), .last_stage(_91[515:515]), .first_stage(_91[514:514]), .start_twiddles(_91[513:513]), .omegas6(_91[512:449]), .omegas5(_91[448:385]), .omegas4(_91[384:321]), .omegas3(_91[320:257]), .omegas2(_91[256:193]), .omegas1(_91[192:129]), .omegas0(_91[128:65]), .addr2(_91[64:53]), .addr1(_91[52:41]), .m(_91[40:29]), .k(_91[28:17]), .j(_91[16:5]), .i(_91[4:1]), .done_(_91[0:0]) );
    assign _1756 = _91[0:0];

    /* aliases */
    assign data_0 = data;
    assign data_2 = data_1;
    assign data_4 = data_3;
    assign data_5 = data_3;
    assign data_6 = data_3;
    assign data_8 = data_7;
    assign data_9 = data_7;
    assign data_10 = data_7;
    assign data_12 = data_11;
    assign data_14 = data_13;
    assign data_16 = data_15;
    assign data_17 = data_15;
    assign data_18 = data_15;
    assign data_20 = data_19;
    assign data_21 = data_19;
    assign data_22 = data_19;
    assign data_24 = data_23;
    assign data_26 = data_25;
    assign data_28 = data_27;
    assign data_29 = data_27;
    assign data_30 = data_27;
    assign data_32 = data_31;
    assign data_33 = data_31;
    assign data_34 = data_31;
    assign data_36 = data_35;
    assign data_38 = data_37;
    assign data_40 = data_39;
    assign data_41 = data_39;
    assign data_42 = data_39;
    assign data_44 = data_43;
    assign data_45 = data_43;
    assign data_46 = data_43;
    assign data_48 = data_47;
    assign data_50 = data_49;
    assign data_52 = data_51;
    assign data_53 = data_51;
    assign data_54 = data_51;
    assign data_56 = data_55;
    assign data_57 = data_55;
    assign data_58 = data_55;
    assign data_60 = data_59;
    assign data_62 = data_61;
    assign data_64 = data_63;
    assign data_65 = data_63;
    assign data_66 = data_63;
    assign data_68 = data_67;
    assign data_69 = data_67;
    assign data_70 = data_67;
    assign data_72 = data_71;
    assign data_74 = data_73;
    assign data_76 = data_75;
    assign data_77 = data_75;
    assign data_78 = data_75;
    assign data_80 = data_79;
    assign data_81 = data_79;
    assign data_82 = data_79;
    assign data_84 = data_83;
    assign data_86 = data_85;
    assign data_88 = data_87;
    assign data_89 = data_87;
    assign data_90 = data_87;
    assign data_92 = data_91;
    assign data_93 = data_91;
    assign data_94 = data_91;

    /* output assignments */
    assign done_ = _1756;
    assign rd_q0 = _1755;
    assign rd_q1 = _1559;
    assign rd_q2 = _1363;
    assign rd_q3 = _1167;
    assign rd_q4 = _971;
    assign rd_q5 = _775;
    assign rd_q6 = _579;
    assign rd_q7 = _383;

endmodule
module dp_39 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1010011101011010110000101010010100001010011101010010100011111111;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0000010100000011100011000110011101011000001110100111010001011001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0001011001000100000110101011001011011010101100111100000011000001;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0100010101011101011101010011001111101010110011010001000101010111;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0101001110010000111001101101001110111101111110001100111010111111;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0010000100011110110101100011101101010010011110100001110000110111;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1100111100000101001110011010010101001111101000110101101001010101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_40 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0110100100111010100111010000000100001110100001110111100100100100;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0000101001101101100000011010111010011001101100111011100011110010;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1111000001010101001011011000111000100001001011011000111001101110;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1111110010010010010101100111111010010010001101101010100101000011;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1111010010000011000001101111100111101101010001110001011010100101;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0101000110110101111111000100110011011110100010011110110011100111;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1100111100101111110001000000111101101011000110000000011001111011;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_41 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0000101110000011010000000101110111010110101101011011110001111001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0011000101111100111000111101000110001100011110101101101000010101;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0011110101010010010000101110111110001011011110110110010010111001;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1011011110011011001100001001011100001010101001010000110000111110;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1110000101110100011000000100000100110100000010000010100100010011;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0110001110111000011110101101110010111010001011110110000001100110;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0010101001001000011111010001011101101011111100000111111100100010;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_42 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0011010001111101110000011100111011011100101110111110011010110111;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1100111011101001011000100111001111100100011101111011111100110001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1000001100110001010001100111100100111111101111100001101111000010;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1110110001001100010000000100110100011011001000100111011100111100;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1010000100011001011000111011101000110101001001011100101011001101;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0100101000100011110001011011000110000100001011000100111010001100;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1111010101100100110100010100000111100100100010001001111010100001;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_43 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0101001100010110000011001010111000110111110101100110100001101001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1001011100000010111011001000011010100101001101110010010110010001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0010000101110010001101000110101010000001001100100101001010100011;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0101011101100100000001000010111010001001011100010100101100010001;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0100011111101001000011110000001000111010101011110101010100100101;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1100101000011000110011110101000000110000010010010011001010001001;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1101101000101011101011101011110001010010100001010000110110101000;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_44 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1100101001000111101011100101000000010101001011001001001000010000;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1111000101010111111011100011110110011011001000100001010100111100;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1010110111100110011000100010011100011010000000110010101000000111;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1010101100000000110010110011010110110001111111010100000010011110;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1010010010110110101001100110111001101110101111010101100100111011;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0100000110110111010100110011011100010101000101100000000101100101;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0101010110001110111110001100010010001010101000010011001111000110;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_45 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1010110011011110000101100010011011111000011011010100011101111000;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0010010101011011011101111010100000000101101000001111000010101010;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1100100001111110110101001111111111010110101111011001101111010010;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0001001110001100011011101101100001010001011001101011101111110100;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0001011011010010100001100000100011010110001111011101101100101001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0001001001101101010000000010001001100101110100000011001111101011;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1010110100011111111111000101110001001001010010010001100001101110;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_46 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1011001000101001010111110011011100011011011110110011111100100000;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1010110110000010101001010101000001011010100011111110110111110010;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0001011001101101101010101011100111100000011110111101111110000010;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1110010101011110011111101111010110001000101101111011011011011101;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1011101010010111101011111110001110001101011101010101011110101010;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1110001001111001110100001100100010011000100011111011110111011010;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1010110100110000000000001100000000101001001101000000111111010000;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module parallel_cores_4 (
    wr_d7,
    wr_d6,
    wr_d5,
    wr_d4,
    wr_d3,
    wr_d2,
    wr_d1,
    wr_d0,
    wr_addr,
    wr_en,
    rd_addr,
    rd_en,
    flip,
    first_4step_pass,
    first_iter,
    start,
    clear,
    clock,
    done_,
    rd_q0,
    rd_q1,
    rd_q2,
    rd_q3,
    rd_q4,
    rd_q5,
    rd_q6,
    rd_q7
);

    input [63:0] wr_d7;
    input [63:0] wr_d6;
    input [63:0] wr_d5;
    input [63:0] wr_d4;
    input [63:0] wr_d3;
    input [63:0] wr_d2;
    input [63:0] wr_d1;
    input [63:0] wr_d0;
    input [11:0] wr_addr;
    input [7:0] wr_en;
    input [11:0] rd_addr;
    input [7:0] rd_en;
    input flip;
    input first_4step_pass;
    input first_iter;
    input start;
    input clear;
    input clock;
    output done_;
    output [63:0] rd_q0;
    output [63:0] rd_q1;
    output [63:0] rd_q2;
    output [63:0] rd_q3;
    output [63:0] rd_q4;
    output [63:0] rd_q5;
    output [63:0] rd_q6;
    output [63:0] rd_q7;

    /* signal declarations */
    wire [11:0] address;
    wire write_enable;
    wire [11:0] address_0;
    wire _374;
    wire read_enable;
    wire _372;
    wire write_enable_0;
    wire _376;
    wire [131:0] _381;
    wire [63:0] _382;
    wire [11:0] _367 = 12'b000000000000;
    wire [11:0] address_1;
    wire _365;
    wire write_enable_1;
    wire [63:0] _279;
    wire [63:0] _278;
    wire [63:0] _280;
    wire [63:0] _276;
    wire [63:0] _275;
    wire [63:0] q1;
    wire [63:0] _281;
    wire [11:0] address_2;
    wire write_enable_2 = 1'b0;
    wire _266;
    wire read_enable_0;
    wire [11:0] address_3;
    wire _262;
    wire read_enable_1;
    wire _260;
    wire write_enable_3;
    wire _264;
    wire [131:0] _271;
    wire [63:0] _272;
    wire [63:0] data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_0;
    wire [11:0] _254 = 12'b000000000000;
    wire _252;
    wire _251;
    wire _250;
    wire _249;
    wire _248;
    wire _247;
    wire _246;
    wire _245;
    wire _244;
    wire _243;
    wire _242;
    wire _241;
    wire [11:0] _253;
    wire [11:0] address_4;
    wire write_enable_4 = 1'b0;
    wire _238;
    wire read_enable_2;
    wire [63:0] data_1;
    wire [63:0] data_2;
    wire _235;
    wire _234;
    wire _233;
    wire _232;
    wire _231;
    wire _230;
    wire _229;
    wire _228;
    wire _227;
    wire _226;
    wire _225;
    wire _224;
    wire [11:0] _236;
    wire [11:0] address_5;
    wire _221;
    wire read_enable_3;
    wire _219;
    wire write_enable_5;
    wire _223;
    wire [131:0] _258;
    wire [63:0] _259;
    wire _87 = 1'b0;
    wire _86 = 1'b0;
    wire _89;
    wire _3;
    reg PHASE;
    wire [63:0] _273;
    wire [11:0] address_6;
    wire _211;
    wire read_enable_4;
    wire write_enable_6;
    wire _213;
    wire [11:0] address_7;
    wire _206;
    wire read_enable_5;
    wire _204;
    wire write_enable_7;
    wire _208;
    wire [131:0] _216;
    wire [63:0] _217;
    wire [63:0] _295;
    wire [63:0] data_3;
    wire [63:0] data_4;
    wire [63:0] data_5;
    wire [63:0] data_6;
    wire [11:0] address_8;
    wire _169;
    wire read_enable_6;
    wire _166;
    wire _167;
    wire write_enable_8;
    wire _171;
    wire [11:0] address_9;
    wire _134;
    wire read_enable_7;
    wire _131;
    wire _132;
    wire write_enable_9;
    wire _136;
    wire [131:0] _202;
    wire [63:0] _203;
    wire _98 = 1'b0;
    wire _97 = 1'b0;
    wire _296;
    wire _5;
    reg PHASE_0;
    wire [63:0] q0;
    wire _94 = 1'b0;
    wire _93 = 1'b0;
    reg _96;
    wire [63:0] _274;
    wire [191:0] _294;
    wire [63:0] _297;
    wire [63:0] data_7;
    wire [63:0] data_8;
    wire [63:0] data_9;
    wire [63:0] data_10;
    wire [11:0] address_10;
    wire _361;
    wire _360;
    wire read_enable_8;
    wire _354 = 1'b0;
    wire _353 = 1'b0;
    wire _351 = 1'b0;
    wire _350 = 1'b0;
    wire _348 = 1'b0;
    wire _347 = 1'b0;
    wire _345 = 1'b0;
    wire _344 = 1'b0;
    wire _342 = 1'b0;
    wire _341 = 1'b0;
    wire _339 = 1'b0;
    wire _338 = 1'b0;
    wire _336 = 1'b0;
    wire _335 = 1'b0;
    wire _333 = 1'b0;
    wire _332 = 1'b0;
    wire _330 = 1'b0;
    wire _329 = 1'b0;
    reg _331;
    reg _334;
    reg _337;
    reg _340;
    reg _343;
    reg _346;
    reg _349;
    reg _352;
    reg _355;
    wire _356;
    wire _327 = 1'b0;
    wire _326 = 1'b0;
    wire _324 = 1'b0;
    wire _323 = 1'b0;
    wire _321 = 1'b0;
    wire _320 = 1'b0;
    wire _318 = 1'b0;
    wire _317 = 1'b0;
    wire _315 = 1'b0;
    wire _314 = 1'b0;
    wire _312 = 1'b0;
    wire _311 = 1'b0;
    wire _309 = 1'b0;
    wire _308 = 1'b0;
    wire _306 = 1'b0;
    wire _305 = 1'b0;
    wire _303 = 1'b0;
    wire _302 = 1'b0;
    reg _304;
    reg _307;
    reg _310;
    reg _313;
    reg _316;
    reg _319;
    reg _322;
    reg _325;
    reg _328;
    wire _357;
    wire _358;
    wire write_enable_10;
    wire _363;
    wire [131:0] _370;
    wire [63:0] _371;
    wire _299 = 1'b0;
    wire _298 = 1'b0;
    wire _301;
    wire _7;
    reg PHASE_1;
    wire [63:0] _383;
    wire [11:0] address_11;
    wire write_enable_11;
    wire [11:0] address_12;
    wire _570;
    wire read_enable_9;
    wire _568;
    wire write_enable_12;
    wire _572;
    wire [131:0] _577;
    wire [63:0] _578;
    wire [11:0] _563 = 12'b000000000000;
    wire [11:0] address_13;
    wire _561;
    wire write_enable_13;
    wire [63:0] _486;
    wire [63:0] _485;
    wire [63:0] _487;
    wire [63:0] _483;
    wire [63:0] _482;
    wire [63:0] q1_0;
    wire [63:0] _488;
    wire [11:0] address_14;
    wire write_enable_14 = 1'b0;
    wire _473;
    wire read_enable_10;
    wire [11:0] address_15;
    wire _469;
    wire read_enable_11;
    wire _467;
    wire write_enable_15;
    wire _471;
    wire [131:0] _478;
    wire [63:0] _479;
    wire [63:0] data_11 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_12;
    wire [11:0] _461 = 12'b000000000000;
    wire _459;
    wire _458;
    wire _457;
    wire _456;
    wire _455;
    wire _454;
    wire _453;
    wire _452;
    wire _451;
    wire _450;
    wire _449;
    wire _448;
    wire [11:0] _460;
    wire [11:0] address_16;
    wire write_enable_16 = 1'b0;
    wire _445;
    wire read_enable_12;
    wire [63:0] data_13;
    wire [63:0] data_14;
    wire _442;
    wire _441;
    wire _440;
    wire _439;
    wire _438;
    wire _437;
    wire _436;
    wire _435;
    wire _434;
    wire _433;
    wire _432;
    wire _431;
    wire [11:0] _443;
    wire [11:0] address_17;
    wire _428;
    wire read_enable_13;
    wire _426;
    wire write_enable_17;
    wire _430;
    wire [131:0] _465;
    wire [63:0] _466;
    wire _385 = 1'b0;
    wire _384 = 1'b0;
    wire _387;
    wire _11;
    reg PHASE_2;
    wire [63:0] _480;
    wire [11:0] address_18;
    wire _418;
    wire read_enable_14;
    wire write_enable_18;
    wire _420;
    wire [11:0] address_19;
    wire _413;
    wire read_enable_15;
    wire _411;
    wire write_enable_19;
    wire _415;
    wire [131:0] _423;
    wire [63:0] _424;
    wire [63:0] _491;
    wire [63:0] data_15;
    wire [63:0] data_16;
    wire [63:0] data_17;
    wire [63:0] data_18;
    wire [11:0] address_20;
    wire _404;
    wire read_enable_16;
    wire _401;
    wire _402;
    wire write_enable_20;
    wire _406;
    wire [11:0] address_21;
    wire _397;
    wire read_enable_17;
    wire _394;
    wire _395;
    wire write_enable_21;
    wire _399;
    wire [131:0] _409;
    wire [63:0] _410;
    wire _392 = 1'b0;
    wire _391 = 1'b0;
    wire _492;
    wire _13;
    reg PHASE_3;
    wire [63:0] q0_0;
    wire _389 = 1'b0;
    wire _388 = 1'b0;
    reg _390;
    wire [63:0] _481;
    wire [191:0] _490;
    wire [63:0] _493;
    wire [63:0] data_19;
    wire [63:0] data_20;
    wire [63:0] data_21;
    wire [63:0] data_22;
    wire [11:0] address_22;
    wire _557;
    wire _556;
    wire read_enable_18;
    wire _550 = 1'b0;
    wire _549 = 1'b0;
    wire _547 = 1'b0;
    wire _546 = 1'b0;
    wire _544 = 1'b0;
    wire _543 = 1'b0;
    wire _541 = 1'b0;
    wire _540 = 1'b0;
    wire _538 = 1'b0;
    wire _537 = 1'b0;
    wire _535 = 1'b0;
    wire _534 = 1'b0;
    wire _532 = 1'b0;
    wire _531 = 1'b0;
    wire _529 = 1'b0;
    wire _528 = 1'b0;
    wire _526 = 1'b0;
    wire _525 = 1'b0;
    reg _527;
    reg _530;
    reg _533;
    reg _536;
    reg _539;
    reg _542;
    reg _545;
    reg _548;
    reg _551;
    wire _552;
    wire _523 = 1'b0;
    wire _522 = 1'b0;
    wire _520 = 1'b0;
    wire _519 = 1'b0;
    wire _517 = 1'b0;
    wire _516 = 1'b0;
    wire _514 = 1'b0;
    wire _513 = 1'b0;
    wire _511 = 1'b0;
    wire _510 = 1'b0;
    wire _508 = 1'b0;
    wire _507 = 1'b0;
    wire _505 = 1'b0;
    wire _504 = 1'b0;
    wire _502 = 1'b0;
    wire _501 = 1'b0;
    wire _499 = 1'b0;
    wire _498 = 1'b0;
    reg _500;
    reg _503;
    reg _506;
    reg _509;
    reg _512;
    reg _515;
    reg _518;
    reg _521;
    reg _524;
    wire _553;
    wire _554;
    wire write_enable_22;
    wire _559;
    wire [131:0] _566;
    wire [63:0] _567;
    wire _495 = 1'b0;
    wire _494 = 1'b0;
    wire _497;
    wire _15;
    reg PHASE_4;
    wire [63:0] _579;
    wire [11:0] address_23;
    wire write_enable_23;
    wire [11:0] address_24;
    wire _766;
    wire read_enable_19;
    wire _764;
    wire write_enable_24;
    wire _768;
    wire [131:0] _773;
    wire [63:0] _774;
    wire [11:0] _759 = 12'b000000000000;
    wire [11:0] address_25;
    wire _757;
    wire write_enable_25;
    wire [63:0] _682;
    wire [63:0] _681;
    wire [63:0] _683;
    wire [63:0] _679;
    wire [63:0] _678;
    wire [63:0] q1_1;
    wire [63:0] _684;
    wire [11:0] address_26;
    wire write_enable_26 = 1'b0;
    wire _669;
    wire read_enable_20;
    wire [11:0] address_27;
    wire _665;
    wire read_enable_21;
    wire _663;
    wire write_enable_27;
    wire _667;
    wire [131:0] _674;
    wire [63:0] _675;
    wire [63:0] data_23 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_24;
    wire [11:0] _657 = 12'b000000000000;
    wire _655;
    wire _654;
    wire _653;
    wire _652;
    wire _651;
    wire _650;
    wire _649;
    wire _648;
    wire _647;
    wire _646;
    wire _645;
    wire _644;
    wire [11:0] _656;
    wire [11:0] address_28;
    wire write_enable_28 = 1'b0;
    wire _641;
    wire read_enable_22;
    wire [63:0] data_25;
    wire [63:0] data_26;
    wire _638;
    wire _637;
    wire _636;
    wire _635;
    wire _634;
    wire _633;
    wire _632;
    wire _631;
    wire _630;
    wire _629;
    wire _628;
    wire _627;
    wire [11:0] _639;
    wire [11:0] address_29;
    wire _624;
    wire read_enable_23;
    wire _622;
    wire write_enable_29;
    wire _626;
    wire [131:0] _661;
    wire [63:0] _662;
    wire _581 = 1'b0;
    wire _580 = 1'b0;
    wire _583;
    wire _19;
    reg PHASE_5;
    wire [63:0] _676;
    wire [11:0] address_30;
    wire _614;
    wire read_enable_24;
    wire write_enable_30;
    wire _616;
    wire [11:0] address_31;
    wire _609;
    wire read_enable_25;
    wire _607;
    wire write_enable_31;
    wire _611;
    wire [131:0] _619;
    wire [63:0] _620;
    wire [63:0] _687;
    wire [63:0] data_27;
    wire [63:0] data_28;
    wire [63:0] data_29;
    wire [63:0] data_30;
    wire [11:0] address_32;
    wire _600;
    wire read_enable_26;
    wire _597;
    wire _598;
    wire write_enable_32;
    wire _602;
    wire [11:0] address_33;
    wire _593;
    wire read_enable_27;
    wire _590;
    wire _591;
    wire write_enable_33;
    wire _595;
    wire [131:0] _605;
    wire [63:0] _606;
    wire _588 = 1'b0;
    wire _587 = 1'b0;
    wire _688;
    wire _21;
    reg PHASE_6;
    wire [63:0] q0_1;
    wire _585 = 1'b0;
    wire _584 = 1'b0;
    reg _586;
    wire [63:0] _677;
    wire [191:0] _686;
    wire [63:0] _689;
    wire [63:0] data_31;
    wire [63:0] data_32;
    wire [63:0] data_33;
    wire [63:0] data_34;
    wire [11:0] address_34;
    wire _753;
    wire _752;
    wire read_enable_28;
    wire _746 = 1'b0;
    wire _745 = 1'b0;
    wire _743 = 1'b0;
    wire _742 = 1'b0;
    wire _740 = 1'b0;
    wire _739 = 1'b0;
    wire _737 = 1'b0;
    wire _736 = 1'b0;
    wire _734 = 1'b0;
    wire _733 = 1'b0;
    wire _731 = 1'b0;
    wire _730 = 1'b0;
    wire _728 = 1'b0;
    wire _727 = 1'b0;
    wire _725 = 1'b0;
    wire _724 = 1'b0;
    wire _722 = 1'b0;
    wire _721 = 1'b0;
    reg _723;
    reg _726;
    reg _729;
    reg _732;
    reg _735;
    reg _738;
    reg _741;
    reg _744;
    reg _747;
    wire _748;
    wire _719 = 1'b0;
    wire _718 = 1'b0;
    wire _716 = 1'b0;
    wire _715 = 1'b0;
    wire _713 = 1'b0;
    wire _712 = 1'b0;
    wire _710 = 1'b0;
    wire _709 = 1'b0;
    wire _707 = 1'b0;
    wire _706 = 1'b0;
    wire _704 = 1'b0;
    wire _703 = 1'b0;
    wire _701 = 1'b0;
    wire _700 = 1'b0;
    wire _698 = 1'b0;
    wire _697 = 1'b0;
    wire _695 = 1'b0;
    wire _694 = 1'b0;
    reg _696;
    reg _699;
    reg _702;
    reg _705;
    reg _708;
    reg _711;
    reg _714;
    reg _717;
    reg _720;
    wire _749;
    wire _750;
    wire write_enable_34;
    wire _755;
    wire [131:0] _762;
    wire [63:0] _763;
    wire _691 = 1'b0;
    wire _690 = 1'b0;
    wire _693;
    wire _23;
    reg PHASE_7;
    wire [63:0] _775;
    wire [11:0] address_35;
    wire write_enable_35;
    wire [11:0] address_36;
    wire _962;
    wire read_enable_29;
    wire _960;
    wire write_enable_36;
    wire _964;
    wire [131:0] _969;
    wire [63:0] _970;
    wire [11:0] _955 = 12'b000000000000;
    wire [11:0] address_37;
    wire _953;
    wire write_enable_37;
    wire [63:0] _878;
    wire [63:0] _877;
    wire [63:0] _879;
    wire [63:0] _875;
    wire [63:0] _874;
    wire [63:0] q1_2;
    wire [63:0] _880;
    wire [11:0] address_38;
    wire write_enable_38 = 1'b0;
    wire _865;
    wire read_enable_30;
    wire [11:0] address_39;
    wire _861;
    wire read_enable_31;
    wire _859;
    wire write_enable_39;
    wire _863;
    wire [131:0] _870;
    wire [63:0] _871;
    wire [63:0] data_35 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_36;
    wire [11:0] _853 = 12'b000000000000;
    wire _851;
    wire _850;
    wire _849;
    wire _848;
    wire _847;
    wire _846;
    wire _845;
    wire _844;
    wire _843;
    wire _842;
    wire _841;
    wire _840;
    wire [11:0] _852;
    wire [11:0] address_40;
    wire write_enable_40 = 1'b0;
    wire _837;
    wire read_enable_32;
    wire [63:0] data_37;
    wire [63:0] data_38;
    wire _834;
    wire _833;
    wire _832;
    wire _831;
    wire _830;
    wire _829;
    wire _828;
    wire _827;
    wire _826;
    wire _825;
    wire _824;
    wire _823;
    wire [11:0] _835;
    wire [11:0] address_41;
    wire _820;
    wire read_enable_33;
    wire _818;
    wire write_enable_41;
    wire _822;
    wire [131:0] _857;
    wire [63:0] _858;
    wire _777 = 1'b0;
    wire _776 = 1'b0;
    wire _779;
    wire _27;
    reg PHASE_8;
    wire [63:0] _872;
    wire [11:0] address_42;
    wire _810;
    wire read_enable_34;
    wire write_enable_42;
    wire _812;
    wire [11:0] address_43;
    wire _805;
    wire read_enable_35;
    wire _803;
    wire write_enable_43;
    wire _807;
    wire [131:0] _815;
    wire [63:0] _816;
    wire [63:0] _883;
    wire [63:0] data_39;
    wire [63:0] data_40;
    wire [63:0] data_41;
    wire [63:0] data_42;
    wire [11:0] address_44;
    wire _796;
    wire read_enable_36;
    wire _793;
    wire _794;
    wire write_enable_44;
    wire _798;
    wire [11:0] address_45;
    wire _789;
    wire read_enable_37;
    wire _786;
    wire _787;
    wire write_enable_45;
    wire _791;
    wire [131:0] _801;
    wire [63:0] _802;
    wire _784 = 1'b0;
    wire _783 = 1'b0;
    wire _884;
    wire _29;
    reg PHASE_9;
    wire [63:0] q0_2;
    wire _781 = 1'b0;
    wire _780 = 1'b0;
    reg _782;
    wire [63:0] _873;
    wire [191:0] _882;
    wire [63:0] _885;
    wire [63:0] data_43;
    wire [63:0] data_44;
    wire [63:0] data_45;
    wire [63:0] data_46;
    wire [11:0] address_46;
    wire _949;
    wire _948;
    wire read_enable_38;
    wire _942 = 1'b0;
    wire _941 = 1'b0;
    wire _939 = 1'b0;
    wire _938 = 1'b0;
    wire _936 = 1'b0;
    wire _935 = 1'b0;
    wire _933 = 1'b0;
    wire _932 = 1'b0;
    wire _930 = 1'b0;
    wire _929 = 1'b0;
    wire _927 = 1'b0;
    wire _926 = 1'b0;
    wire _924 = 1'b0;
    wire _923 = 1'b0;
    wire _921 = 1'b0;
    wire _920 = 1'b0;
    wire _918 = 1'b0;
    wire _917 = 1'b0;
    reg _919;
    reg _922;
    reg _925;
    reg _928;
    reg _931;
    reg _934;
    reg _937;
    reg _940;
    reg _943;
    wire _944;
    wire _915 = 1'b0;
    wire _914 = 1'b0;
    wire _912 = 1'b0;
    wire _911 = 1'b0;
    wire _909 = 1'b0;
    wire _908 = 1'b0;
    wire _906 = 1'b0;
    wire _905 = 1'b0;
    wire _903 = 1'b0;
    wire _902 = 1'b0;
    wire _900 = 1'b0;
    wire _899 = 1'b0;
    wire _897 = 1'b0;
    wire _896 = 1'b0;
    wire _894 = 1'b0;
    wire _893 = 1'b0;
    wire _891 = 1'b0;
    wire _890 = 1'b0;
    reg _892;
    reg _895;
    reg _898;
    reg _901;
    reg _904;
    reg _907;
    reg _910;
    reg _913;
    reg _916;
    wire _945;
    wire _946;
    wire write_enable_46;
    wire _951;
    wire [131:0] _958;
    wire [63:0] _959;
    wire _887 = 1'b0;
    wire _886 = 1'b0;
    wire _889;
    wire _31;
    reg PHASE_10;
    wire [63:0] _971;
    wire [11:0] address_47;
    wire write_enable_47;
    wire [11:0] address_48;
    wire _1158;
    wire read_enable_39;
    wire _1156;
    wire write_enable_48;
    wire _1160;
    wire [131:0] _1165;
    wire [63:0] _1166;
    wire [11:0] _1151 = 12'b000000000000;
    wire [11:0] address_49;
    wire _1149;
    wire write_enable_49;
    wire [63:0] _1074;
    wire [63:0] _1073;
    wire [63:0] _1075;
    wire [63:0] _1071;
    wire [63:0] _1070;
    wire [63:0] q1_3;
    wire [63:0] _1076;
    wire [11:0] address_50;
    wire write_enable_50 = 1'b0;
    wire _1061;
    wire read_enable_40;
    wire [11:0] address_51;
    wire _1057;
    wire read_enable_41;
    wire _1055;
    wire write_enable_51;
    wire _1059;
    wire [131:0] _1066;
    wire [63:0] _1067;
    wire [63:0] data_47 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_48;
    wire [11:0] _1049 = 12'b000000000000;
    wire _1047;
    wire _1046;
    wire _1045;
    wire _1044;
    wire _1043;
    wire _1042;
    wire _1041;
    wire _1040;
    wire _1039;
    wire _1038;
    wire _1037;
    wire _1036;
    wire [11:0] _1048;
    wire [11:0] address_52;
    wire write_enable_52 = 1'b0;
    wire _1033;
    wire read_enable_42;
    wire [63:0] data_49;
    wire [63:0] data_50;
    wire _1030;
    wire _1029;
    wire _1028;
    wire _1027;
    wire _1026;
    wire _1025;
    wire _1024;
    wire _1023;
    wire _1022;
    wire _1021;
    wire _1020;
    wire _1019;
    wire [11:0] _1031;
    wire [11:0] address_53;
    wire _1016;
    wire read_enable_43;
    wire _1014;
    wire write_enable_53;
    wire _1018;
    wire [131:0] _1053;
    wire [63:0] _1054;
    wire _973 = 1'b0;
    wire _972 = 1'b0;
    wire _975;
    wire _35;
    reg PHASE_11;
    wire [63:0] _1068;
    wire [11:0] address_54;
    wire _1006;
    wire read_enable_44;
    wire write_enable_54;
    wire _1008;
    wire [11:0] address_55;
    wire _1001;
    wire read_enable_45;
    wire _999;
    wire write_enable_55;
    wire _1003;
    wire [131:0] _1011;
    wire [63:0] _1012;
    wire [63:0] _1079;
    wire [63:0] data_51;
    wire [63:0] data_52;
    wire [63:0] data_53;
    wire [63:0] data_54;
    wire [11:0] address_56;
    wire _992;
    wire read_enable_46;
    wire _989;
    wire _990;
    wire write_enable_56;
    wire _994;
    wire [11:0] address_57;
    wire _985;
    wire read_enable_47;
    wire _982;
    wire _983;
    wire write_enable_57;
    wire _987;
    wire [131:0] _997;
    wire [63:0] _998;
    wire _980 = 1'b0;
    wire _979 = 1'b0;
    wire _1080;
    wire _37;
    reg PHASE_12;
    wire [63:0] q0_3;
    wire _977 = 1'b0;
    wire _976 = 1'b0;
    reg _978;
    wire [63:0] _1069;
    wire [191:0] _1078;
    wire [63:0] _1081;
    wire [63:0] data_55;
    wire [63:0] data_56;
    wire [63:0] data_57;
    wire [63:0] data_58;
    wire [11:0] address_58;
    wire _1145;
    wire _1144;
    wire read_enable_48;
    wire _1138 = 1'b0;
    wire _1137 = 1'b0;
    wire _1135 = 1'b0;
    wire _1134 = 1'b0;
    wire _1132 = 1'b0;
    wire _1131 = 1'b0;
    wire _1129 = 1'b0;
    wire _1128 = 1'b0;
    wire _1126 = 1'b0;
    wire _1125 = 1'b0;
    wire _1123 = 1'b0;
    wire _1122 = 1'b0;
    wire _1120 = 1'b0;
    wire _1119 = 1'b0;
    wire _1117 = 1'b0;
    wire _1116 = 1'b0;
    wire _1114 = 1'b0;
    wire _1113 = 1'b0;
    reg _1115;
    reg _1118;
    reg _1121;
    reg _1124;
    reg _1127;
    reg _1130;
    reg _1133;
    reg _1136;
    reg _1139;
    wire _1140;
    wire _1111 = 1'b0;
    wire _1110 = 1'b0;
    wire _1108 = 1'b0;
    wire _1107 = 1'b0;
    wire _1105 = 1'b0;
    wire _1104 = 1'b0;
    wire _1102 = 1'b0;
    wire _1101 = 1'b0;
    wire _1099 = 1'b0;
    wire _1098 = 1'b0;
    wire _1096 = 1'b0;
    wire _1095 = 1'b0;
    wire _1093 = 1'b0;
    wire _1092 = 1'b0;
    wire _1090 = 1'b0;
    wire _1089 = 1'b0;
    wire _1087 = 1'b0;
    wire _1086 = 1'b0;
    reg _1088;
    reg _1091;
    reg _1094;
    reg _1097;
    reg _1100;
    reg _1103;
    reg _1106;
    reg _1109;
    reg _1112;
    wire _1141;
    wire _1142;
    wire write_enable_58;
    wire _1147;
    wire [131:0] _1154;
    wire [63:0] _1155;
    wire _1083 = 1'b0;
    wire _1082 = 1'b0;
    wire _1085;
    wire _39;
    reg PHASE_13;
    wire [63:0] _1167;
    wire [11:0] address_59;
    wire write_enable_59;
    wire [11:0] address_60;
    wire _1354;
    wire read_enable_49;
    wire _1352;
    wire write_enable_60;
    wire _1356;
    wire [131:0] _1361;
    wire [63:0] _1362;
    wire [11:0] _1347 = 12'b000000000000;
    wire [11:0] address_61;
    wire _1345;
    wire write_enable_61;
    wire [63:0] _1270;
    wire [63:0] _1269;
    wire [63:0] _1271;
    wire [63:0] _1267;
    wire [63:0] _1266;
    wire [63:0] q1_4;
    wire [63:0] _1272;
    wire [11:0] address_62;
    wire write_enable_62 = 1'b0;
    wire _1257;
    wire read_enable_50;
    wire [11:0] address_63;
    wire _1253;
    wire read_enable_51;
    wire _1251;
    wire write_enable_63;
    wire _1255;
    wire [131:0] _1262;
    wire [63:0] _1263;
    wire [63:0] data_59 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_60;
    wire [11:0] _1245 = 12'b000000000000;
    wire _1243;
    wire _1242;
    wire _1241;
    wire _1240;
    wire _1239;
    wire _1238;
    wire _1237;
    wire _1236;
    wire _1235;
    wire _1234;
    wire _1233;
    wire _1232;
    wire [11:0] _1244;
    wire [11:0] address_64;
    wire write_enable_64 = 1'b0;
    wire _1229;
    wire read_enable_52;
    wire [63:0] data_61;
    wire [63:0] data_62;
    wire _1226;
    wire _1225;
    wire _1224;
    wire _1223;
    wire _1222;
    wire _1221;
    wire _1220;
    wire _1219;
    wire _1218;
    wire _1217;
    wire _1216;
    wire _1215;
    wire [11:0] _1227;
    wire [11:0] address_65;
    wire _1212;
    wire read_enable_53;
    wire _1210;
    wire write_enable_65;
    wire _1214;
    wire [131:0] _1249;
    wire [63:0] _1250;
    wire _1169 = 1'b0;
    wire _1168 = 1'b0;
    wire _1171;
    wire _43;
    reg PHASE_14;
    wire [63:0] _1264;
    wire [11:0] address_66;
    wire _1202;
    wire read_enable_54;
    wire write_enable_66;
    wire _1204;
    wire [11:0] address_67;
    wire _1197;
    wire read_enable_55;
    wire _1195;
    wire write_enable_67;
    wire _1199;
    wire [131:0] _1207;
    wire [63:0] _1208;
    wire [63:0] _1275;
    wire [63:0] data_63;
    wire [63:0] data_64;
    wire [63:0] data_65;
    wire [63:0] data_66;
    wire [11:0] address_68;
    wire _1188;
    wire read_enable_56;
    wire _1185;
    wire _1186;
    wire write_enable_68;
    wire _1190;
    wire [11:0] address_69;
    wire _1181;
    wire read_enable_57;
    wire _1178;
    wire _1179;
    wire write_enable_69;
    wire _1183;
    wire [131:0] _1193;
    wire [63:0] _1194;
    wire _1176 = 1'b0;
    wire _1175 = 1'b0;
    wire _1276;
    wire _45;
    reg PHASE_15;
    wire [63:0] q0_4;
    wire _1173 = 1'b0;
    wire _1172 = 1'b0;
    reg _1174;
    wire [63:0] _1265;
    wire [191:0] _1274;
    wire [63:0] _1277;
    wire [63:0] data_67;
    wire [63:0] data_68;
    wire [63:0] data_69;
    wire [63:0] data_70;
    wire [11:0] address_70;
    wire _1341;
    wire _1340;
    wire read_enable_58;
    wire _1334 = 1'b0;
    wire _1333 = 1'b0;
    wire _1331 = 1'b0;
    wire _1330 = 1'b0;
    wire _1328 = 1'b0;
    wire _1327 = 1'b0;
    wire _1325 = 1'b0;
    wire _1324 = 1'b0;
    wire _1322 = 1'b0;
    wire _1321 = 1'b0;
    wire _1319 = 1'b0;
    wire _1318 = 1'b0;
    wire _1316 = 1'b0;
    wire _1315 = 1'b0;
    wire _1313 = 1'b0;
    wire _1312 = 1'b0;
    wire _1310 = 1'b0;
    wire _1309 = 1'b0;
    reg _1311;
    reg _1314;
    reg _1317;
    reg _1320;
    reg _1323;
    reg _1326;
    reg _1329;
    reg _1332;
    reg _1335;
    wire _1336;
    wire _1307 = 1'b0;
    wire _1306 = 1'b0;
    wire _1304 = 1'b0;
    wire _1303 = 1'b0;
    wire _1301 = 1'b0;
    wire _1300 = 1'b0;
    wire _1298 = 1'b0;
    wire _1297 = 1'b0;
    wire _1295 = 1'b0;
    wire _1294 = 1'b0;
    wire _1292 = 1'b0;
    wire _1291 = 1'b0;
    wire _1289 = 1'b0;
    wire _1288 = 1'b0;
    wire _1286 = 1'b0;
    wire _1285 = 1'b0;
    wire _1283 = 1'b0;
    wire _1282 = 1'b0;
    reg _1284;
    reg _1287;
    reg _1290;
    reg _1293;
    reg _1296;
    reg _1299;
    reg _1302;
    reg _1305;
    reg _1308;
    wire _1337;
    wire _1338;
    wire write_enable_70;
    wire _1343;
    wire [131:0] _1350;
    wire [63:0] _1351;
    wire _1279 = 1'b0;
    wire _1278 = 1'b0;
    wire _1281;
    wire _47;
    reg PHASE_16;
    wire [63:0] _1363;
    wire [11:0] address_71;
    wire write_enable_71;
    wire [11:0] address_72;
    wire _1550;
    wire read_enable_59;
    wire _1548;
    wire write_enable_72;
    wire _1552;
    wire [131:0] _1557;
    wire [63:0] _1558;
    wire [11:0] _1543 = 12'b000000000000;
    wire [11:0] address_73;
    wire _1541;
    wire write_enable_73;
    wire [63:0] _1466;
    wire [63:0] _1465;
    wire [63:0] _1467;
    wire [63:0] _1463;
    wire [63:0] _1462;
    wire [63:0] q1_5;
    wire [63:0] _1468;
    wire [11:0] address_74;
    wire write_enable_74 = 1'b0;
    wire _1453;
    wire read_enable_60;
    wire [11:0] address_75;
    wire _1449;
    wire read_enable_61;
    wire _1447;
    wire write_enable_75;
    wire _1451;
    wire [131:0] _1458;
    wire [63:0] _1459;
    wire [63:0] data_71 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_72;
    wire [11:0] _1441 = 12'b000000000000;
    wire _1439;
    wire _1438;
    wire _1437;
    wire _1436;
    wire _1435;
    wire _1434;
    wire _1433;
    wire _1432;
    wire _1431;
    wire _1430;
    wire _1429;
    wire _1428;
    wire [11:0] _1440;
    wire [11:0] address_76;
    wire write_enable_76 = 1'b0;
    wire _1425;
    wire read_enable_62;
    wire [63:0] data_73;
    wire [63:0] data_74;
    wire _1422;
    wire _1421;
    wire _1420;
    wire _1419;
    wire _1418;
    wire _1417;
    wire _1416;
    wire _1415;
    wire _1414;
    wire _1413;
    wire _1412;
    wire _1411;
    wire [11:0] _1423;
    wire [11:0] address_77;
    wire _1408;
    wire read_enable_63;
    wire _1406;
    wire write_enable_77;
    wire _1410;
    wire [131:0] _1445;
    wire [63:0] _1446;
    wire _1365 = 1'b0;
    wire _1364 = 1'b0;
    wire _1367;
    wire _51;
    reg PHASE_17;
    wire [63:0] _1460;
    wire [11:0] address_78;
    wire _1398;
    wire read_enable_64;
    wire write_enable_78;
    wire _1400;
    wire [11:0] address_79;
    wire _1393;
    wire read_enable_65;
    wire _1391;
    wire write_enable_79;
    wire _1395;
    wire [131:0] _1403;
    wire [63:0] _1404;
    wire [63:0] _1471;
    wire [63:0] data_75;
    wire [63:0] data_76;
    wire [63:0] data_77;
    wire [63:0] data_78;
    wire [11:0] address_80;
    wire _1384;
    wire read_enable_66;
    wire _1381;
    wire _1382;
    wire write_enable_80;
    wire _1386;
    wire [11:0] address_81;
    wire _1377;
    wire read_enable_67;
    wire _1374;
    wire _1375;
    wire write_enable_81;
    wire _1379;
    wire [131:0] _1389;
    wire [63:0] _1390;
    wire _1372 = 1'b0;
    wire _1371 = 1'b0;
    wire _1472;
    wire _53;
    reg PHASE_18;
    wire [63:0] q0_5;
    wire _1369 = 1'b0;
    wire _1368 = 1'b0;
    reg _1370;
    wire [63:0] _1461;
    wire [191:0] _1470;
    wire [63:0] _1473;
    wire [63:0] data_79;
    wire [63:0] data_80;
    wire [63:0] data_81;
    wire [63:0] data_82;
    wire [11:0] address_82;
    wire _1537;
    wire _1536;
    wire read_enable_68;
    wire _1530 = 1'b0;
    wire _1529 = 1'b0;
    wire _1527 = 1'b0;
    wire _1526 = 1'b0;
    wire _1524 = 1'b0;
    wire _1523 = 1'b0;
    wire _1521 = 1'b0;
    wire _1520 = 1'b0;
    wire _1518 = 1'b0;
    wire _1517 = 1'b0;
    wire _1515 = 1'b0;
    wire _1514 = 1'b0;
    wire _1512 = 1'b0;
    wire _1511 = 1'b0;
    wire _1509 = 1'b0;
    wire _1508 = 1'b0;
    wire _1506 = 1'b0;
    wire _1505 = 1'b0;
    reg _1507;
    reg _1510;
    reg _1513;
    reg _1516;
    reg _1519;
    reg _1522;
    reg _1525;
    reg _1528;
    reg _1531;
    wire _1532;
    wire _1503 = 1'b0;
    wire _1502 = 1'b0;
    wire _1500 = 1'b0;
    wire _1499 = 1'b0;
    wire _1497 = 1'b0;
    wire _1496 = 1'b0;
    wire _1494 = 1'b0;
    wire _1493 = 1'b0;
    wire _1491 = 1'b0;
    wire _1490 = 1'b0;
    wire _1488 = 1'b0;
    wire _1487 = 1'b0;
    wire _1485 = 1'b0;
    wire _1484 = 1'b0;
    wire _1482 = 1'b0;
    wire _1481 = 1'b0;
    wire _1479 = 1'b0;
    wire _1478 = 1'b0;
    reg _1480;
    reg _1483;
    reg _1486;
    reg _1489;
    reg _1492;
    reg _1495;
    reg _1498;
    reg _1501;
    reg _1504;
    wire _1533;
    wire _1534;
    wire write_enable_82;
    wire _1539;
    wire [131:0] _1546;
    wire [63:0] _1547;
    wire _1475 = 1'b0;
    wire _1474 = 1'b0;
    wire _1477;
    wire _55;
    reg PHASE_19;
    wire [63:0] _1559;
    wire [11:0] address_83;
    wire write_enable_83;
    wire [11:0] address_84;
    wire _1746;
    wire read_enable_69;
    wire _1744;
    wire write_enable_84;
    wire _1748;
    wire [131:0] _1753;
    wire [63:0] _1754;
    wire [11:0] _1739 = 12'b000000000000;
    wire [11:0] address_85;
    wire _1737;
    wire write_enable_85;
    wire [3:0] _292;
    wire _291;
    wire _289;
    wire [63:0] _288;
    wire [63:0] _287;
    wire [63:0] _286;
    wire [63:0] _285;
    wire [63:0] _284;
    wire [63:0] _283;
    wire [63:0] _282;
    wire [63:0] _1662;
    wire [63:0] _1661;
    wire [63:0] _1663;
    wire [63:0] _1659;
    wire [63:0] _1658;
    wire [63:0] q1_6;
    wire [63:0] _1664;
    wire [11:0] address_86;
    wire write_enable_86 = 1'b0;
    wire _1649;
    wire read_enable_70;
    wire [11:0] address_87;
    wire _1645;
    wire read_enable_71;
    wire _1643;
    wire write_enable_87;
    wire _1647;
    wire [131:0] _1654;
    wire [63:0] _1655;
    wire [63:0] data_83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_84;
    wire [11:0] _1637 = 12'b000000000000;
    wire _1635;
    wire _1634;
    wire _1633;
    wire _1632;
    wire _1631;
    wire _1630;
    wire _1629;
    wire _1628;
    wire _1627;
    wire _1626;
    wire _1625;
    wire _1624;
    wire [11:0] _1636;
    wire [11:0] address_88;
    wire write_enable_88 = 1'b0;
    wire _1621;
    wire read_enable_72;
    wire [63:0] data_85;
    wire [63:0] data_86;
    wire [11:0] _60;
    wire _1618;
    wire _1617;
    wire _1616;
    wire _1615;
    wire _1614;
    wire _1613;
    wire _1612;
    wire _1611;
    wire _1610;
    wire _1609;
    wire _1608;
    wire _1607;
    wire [11:0] _1619;
    wire [11:0] address_89;
    wire _1604;
    wire read_enable_73;
    wire [7:0] _62;
    wire _1602;
    wire write_enable_89;
    wire _1606;
    wire [131:0] _1641;
    wire [63:0] _1642;
    wire _1561 = 1'b0;
    wire _1560 = 1'b0;
    wire _1563;
    wire _63;
    reg PHASE_20;
    wire [63:0] _1656;
    wire [11:0] address_90;
    wire _1594;
    wire read_enable_74;
    wire write_enable_90;
    wire _1596;
    wire [11:0] address_91;
    wire _1589;
    wire read_enable_75;
    wire _1587;
    wire write_enable_91;
    wire _1591;
    wire [131:0] _1599;
    wire [63:0] _1600;
    wire [63:0] _1667;
    wire [63:0] data_87;
    wire [63:0] data_88;
    wire [63:0] data_89;
    wire [63:0] data_90;
    wire [11:0] _198 = 12'b000000000000;
    wire [11:0] _197 = 12'b000000000000;
    wire [11:0] _195 = 12'b000000000000;
    wire [11:0] _194 = 12'b000000000000;
    wire [11:0] _192 = 12'b000000000000;
    wire [11:0] _191 = 12'b000000000000;
    wire [11:0] _189 = 12'b000000000000;
    wire [11:0] _188 = 12'b000000000000;
    wire [11:0] _186 = 12'b000000000000;
    wire [11:0] _185 = 12'b000000000000;
    wire [11:0] _183 = 12'b000000000000;
    wire [11:0] _182 = 12'b000000000000;
    wire [11:0] _180 = 12'b000000000000;
    wire [11:0] _179 = 12'b000000000000;
    wire [11:0] _177 = 12'b000000000000;
    wire [11:0] _176 = 12'b000000000000;
    wire [11:0] _174 = 12'b000000000000;
    wire [11:0] _173 = 12'b000000000000;
    reg [11:0] _175;
    reg [11:0] _178;
    reg [11:0] _181;
    reg [11:0] _184;
    reg [11:0] _187;
    reg [11:0] _190;
    reg [11:0] _193;
    reg [11:0] _196;
    reg [11:0] _199;
    wire [11:0] _172;
    wire [11:0] address_92;
    wire _1580;
    wire read_enable_76;
    wire _1577;
    wire _1578;
    wire write_enable_92;
    wire _1582;
    wire [11:0] address_93;
    wire _1573;
    wire read_enable_77;
    wire _1570;
    wire _1571;
    wire write_enable_93;
    wire _1575;
    wire [131:0] _1585;
    wire [63:0] _1586;
    wire _99;
    wire _1568 = 1'b0;
    wire _1567 = 1'b0;
    wire _1668;
    wire _65;
    reg PHASE_21;
    wire [63:0] q0_6;
    wire _1565 = 1'b0;
    wire _1564 = 1'b0;
    wire _92;
    reg _1566;
    wire [63:0] _1657;
    wire [191:0] _1666;
    wire [63:0] _1669;
    wire [63:0] data_91;
    wire [63:0] data_92;
    wire [63:0] data_93;
    wire [63:0] data_94;
    wire [11:0] _163 = 12'b000000000000;
    wire [11:0] _162 = 12'b000000000000;
    wire [11:0] _160 = 12'b000000000000;
    wire [11:0] _159 = 12'b000000000000;
    wire [11:0] _157 = 12'b000000000000;
    wire [11:0] _156 = 12'b000000000000;
    wire [11:0] _154 = 12'b000000000000;
    wire [11:0] _153 = 12'b000000000000;
    wire [11:0] _151 = 12'b000000000000;
    wire [11:0] _150 = 12'b000000000000;
    wire [11:0] _148 = 12'b000000000000;
    wire [11:0] _147 = 12'b000000000000;
    wire [11:0] _145 = 12'b000000000000;
    wire [11:0] _144 = 12'b000000000000;
    wire [11:0] _142 = 12'b000000000000;
    wire [11:0] _141 = 12'b000000000000;
    wire [11:0] _139 = 12'b000000000000;
    wire [11:0] _138 = 12'b000000000000;
    wire [11:0] _137;
    reg [11:0] _140;
    reg [11:0] _143;
    reg [11:0] _146;
    reg [11:0] _149;
    reg [11:0] _152;
    reg [11:0] _155;
    reg [11:0] _158;
    reg [11:0] _161;
    reg [11:0] _164;
    wire [11:0] _68;
    wire [11:0] address_94;
    wire _1733;
    wire [7:0] _70;
    wire _1732;
    wire read_enable_78;
    wire _1726 = 1'b0;
    wire _1725 = 1'b0;
    wire _1723 = 1'b0;
    wire _1722 = 1'b0;
    wire _1720 = 1'b0;
    wire _1719 = 1'b0;
    wire _1717 = 1'b0;
    wire _1716 = 1'b0;
    wire _1714 = 1'b0;
    wire _1713 = 1'b0;
    wire _1711 = 1'b0;
    wire _1710 = 1'b0;
    wire _1708 = 1'b0;
    wire _1707 = 1'b0;
    wire _1705 = 1'b0;
    wire _1704 = 1'b0;
    wire _1702 = 1'b0;
    wire _1701 = 1'b0;
    wire _290;
    reg _1703;
    reg _1706;
    reg _1709;
    reg _1712;
    reg _1715;
    reg _1718;
    reg _1721;
    reg _1724;
    reg _1727;
    wire _1728;
    wire _1699 = 1'b0;
    wire _1698 = 1'b0;
    wire _1696 = 1'b0;
    wire _1695 = 1'b0;
    wire _1693 = 1'b0;
    wire _1692 = 1'b0;
    wire _1690 = 1'b0;
    wire _1689 = 1'b0;
    wire _1687 = 1'b0;
    wire _1686 = 1'b0;
    wire _1684 = 1'b0;
    wire _1683 = 1'b0;
    wire _1681 = 1'b0;
    wire _1680 = 1'b0;
    wire _1678 = 1'b0;
    wire _1677 = 1'b0;
    wire _1675 = 1'b0;
    wire _1674 = 1'b0;
    wire _130;
    reg _1676;
    reg _1679;
    reg _1682;
    reg _1685;
    reg _1688;
    reg _1691;
    reg _1694;
    reg _1697;
    reg _1700;
    wire _1729;
    wire _128 = 1'b0;
    wire _127 = 1'b0;
    wire _125 = 1'b0;
    wire _124 = 1'b0;
    wire _122 = 1'b0;
    wire _121 = 1'b0;
    wire _119 = 1'b0;
    wire _118 = 1'b0;
    wire _116 = 1'b0;
    wire _115 = 1'b0;
    wire _113 = 1'b0;
    wire _112 = 1'b0;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire vdd = 1'b1;
    wire _104 = 1'b0;
    wire _103 = 1'b0;
    wire _102;
    reg _105;
    reg _108;
    reg _111;
    reg _114;
    reg _117;
    reg _120;
    reg _123;
    reg _126;
    reg _129;
    wire _1730;
    wire write_enable_94;
    wire _1735;
    wire gnd = 1'b0;
    wire [131:0] _1742;
    wire [63:0] _1743;
    wire _72;
    wire _1671 = 1'b0;
    wire _1670 = 1'b0;
    wire _1673;
    wire _73;
    reg PHASE_22;
    wire [63:0] _1755;
    wire _76;
    wire _78;
    wire _80;
    wire _82;
    wire _84;
    wire [523:0] _91;
    wire _1756;

    /* logic */
    assign address = _372 ? _199 : _367;
    assign write_enable = _365 & _372;
    assign address_0 = _372 ? _164 : _68;
    assign _374 = ~ _372;
    assign read_enable = _360 & _374;
    assign _372 = ~ PHASE_1;
    assign write_enable_0 = _358 & _372;
    assign _376 = write_enable_0 | read_enable;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_376), .regcea(vdd), .wea(write_enable_0), .addra(address_0), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable), .regceb(vdd), .web(write_enable), .addrb(address), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_381[131:131]), .sbiterrb(_381[130:130]), .doutb(_381[129:66]), .dbiterra(_381[65:65]), .sbiterra(_381[64:64]), .douta(_381[63:0]) );
    assign _382 = _381[63:0];
    assign address_1 = PHASE_1 ? _199 : _367;
    assign _365 = _129 & _328;
    assign write_enable_1 = _365 & PHASE_1;
    assign _279 = _271[129:66];
    assign _278 = _258[129:66];
    assign _280 = PHASE ? _279 : _278;
    assign _276 = _216[129:66];
    assign _275 = _202[129:66];
    assign q1 = PHASE_0 ? _276 : _275;
    assign _281 = _96 ? _280 : q1;
    assign address_2 = _260 ? _254 : _253;
    assign _266 = ~ _260;
    assign read_enable_0 = _102 & _266;
    assign address_3 = _260 ? _60 : _236;
    assign _262 = ~ _260;
    assign read_enable_1 = _102 & _262;
    assign _260 = ~ PHASE;
    assign write_enable_3 = _219 & _260;
    assign _264 = write_enable_3 | read_enable_1;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_0
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_264), .regcea(vdd), .wea(write_enable_3), .addra(address_3), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_0), .regceb(vdd), .web(write_enable_2), .addrb(address_2), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_271[131:131]), .sbiterrb(_271[130:130]), .doutb(_271[129:66]), .dbiterra(_271[65:65]), .sbiterra(_271[64:64]), .douta(_271[63:0]) );
    assign _272 = _271[63:0];
    assign _252 = _172[11:11];
    assign _251 = _172[10:10];
    assign _250 = _172[9:9];
    assign _249 = _172[8:8];
    assign _248 = _172[7:7];
    assign _247 = _172[6:6];
    assign _246 = _172[5:5];
    assign _245 = _172[4:4];
    assign _244 = _172[3:3];
    assign _243 = _172[2:2];
    assign _242 = _172[1:1];
    assign _241 = _172[0:0];
    assign _253 = { _241, _242, _243, _244, _245, _246, _247, _248, _249, _250, _251, _252 };
    assign address_4 = PHASE ? _254 : _253;
    assign _238 = ~ PHASE;
    assign read_enable_2 = _102 & _238;
    assign data_1 = wr_d7;
    assign _235 = _137[11:11];
    assign _234 = _137[10:10];
    assign _233 = _137[9:9];
    assign _232 = _137[8:8];
    assign _231 = _137[7:7];
    assign _230 = _137[6:6];
    assign _229 = _137[5:5];
    assign _228 = _137[4:4];
    assign _227 = _137[3:3];
    assign _226 = _137[2:2];
    assign _225 = _137[1:1];
    assign _224 = _137[0:0];
    assign _236 = { _224, _225, _226, _227, _228, _229, _230, _231, _232, _233, _234, _235 };
    assign address_5 = PHASE ? _60 : _236;
    assign _221 = ~ PHASE;
    assign read_enable_3 = _102 & _221;
    assign _219 = _62[7:7];
    assign write_enable_5 = _219 & PHASE;
    assign _223 = write_enable_5 | read_enable_3;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_1
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_223), .regcea(vdd), .wea(write_enable_5), .addra(address_5), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_2), .regceb(vdd), .web(write_enable_4), .addrb(address_4), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_258[131:131]), .sbiterrb(_258[130:130]), .doutb(_258[129:66]), .dbiterra(_258[65:65]), .sbiterra(_258[64:64]), .douta(_258[63:0]) );
    assign _259 = _258[63:0];
    assign _89 = ~ PHASE;
    assign _3 = _89;
    always @(posedge _84) begin
        if (_82)
            PHASE <= _87;
        else
            if (_72)
                PHASE <= _3;
    end
    assign _273 = PHASE ? _272 : _259;
    assign address_6 = _204 ? _199 : _172;
    assign _211 = ~ _204;
    assign read_enable_4 = _102 & _211;
    assign write_enable_6 = _167 & _204;
    assign _213 = write_enable_6 | read_enable_4;
    assign address_7 = _204 ? _164 : _137;
    assign _206 = ~ _204;
    assign read_enable_5 = _102 & _206;
    assign _204 = ~ PHASE_0;
    assign write_enable_7 = _132 & _204;
    assign _208 = write_enable_7 | read_enable_5;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_2
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_208), .regcea(vdd), .wea(write_enable_7), .addra(address_7), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_213), .regceb(vdd), .web(write_enable_6), .addrb(address_6), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_216[131:131]), .sbiterrb(_216[130:130]), .doutb(_216[129:66]), .dbiterra(_216[65:65]), .sbiterra(_216[64:64]), .douta(_216[63:0]) );
    assign _217 = _216[63:0];
    assign _295 = _294[127:64];
    assign data_3 = _295;
    assign address_8 = PHASE_0 ? _199 : _172;
    assign _169 = ~ PHASE_0;
    assign read_enable_6 = _102 & _169;
    assign _166 = ~ _130;
    assign _167 = _129 & _166;
    assign write_enable_8 = _167 & PHASE_0;
    assign _171 = write_enable_8 | read_enable_6;
    assign address_9 = PHASE_0 ? _164 : _137;
    assign _134 = ~ PHASE_0;
    assign read_enable_7 = _102 & _134;
    assign _131 = ~ _130;
    assign _132 = _129 & _131;
    assign write_enable_9 = _132 & PHASE_0;
    assign _136 = write_enable_9 | read_enable_7;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_3
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_136), .regcea(vdd), .wea(write_enable_9), .addra(address_9), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_171), .regceb(vdd), .web(write_enable_8), .addrb(address_8), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_202[131:131]), .sbiterrb(_202[130:130]), .doutb(_202[129:66]), .dbiterra(_202[65:65]), .sbiterra(_202[64:64]), .douta(_202[63:0]) );
    assign _203 = _202[63:0];
    assign _296 = ~ PHASE_0;
    assign _5 = _296;
    always @(posedge _84) begin
        if (_82)
            PHASE_0 <= _98;
        else
            if (_99)
                PHASE_0 <= _5;
    end
    assign q0 = PHASE_0 ? _217 : _203;
    always @(posedge _84) begin
        if (_82)
            _96 <= _94;
        else
            _96 <= _92;
    end
    assign _274 = _96 ? _273 : q0;
    dp_46
        dp_6
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_274), .d2(_281), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_294[191:128]), .q2(_294[127:64]), .q1(_294[63:0]) );
    assign _297 = _294[63:0];
    assign data_7 = _297;
    assign address_10 = PHASE_1 ? _164 : _68;
    assign _361 = ~ PHASE_1;
    assign _360 = _70[7:7];
    assign read_enable_8 = _360 & _361;
    always @(posedge _84) begin
        if (_82)
            _331 <= _330;
        else
            _331 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _334 <= _333;
        else
            _334 <= _331;
    end
    always @(posedge _84) begin
        if (_82)
            _337 <= _336;
        else
            _337 <= _334;
    end
    always @(posedge _84) begin
        if (_82)
            _340 <= _339;
        else
            _340 <= _337;
    end
    always @(posedge _84) begin
        if (_82)
            _343 <= _342;
        else
            _343 <= _340;
    end
    always @(posedge _84) begin
        if (_82)
            _346 <= _345;
        else
            _346 <= _343;
    end
    always @(posedge _84) begin
        if (_82)
            _349 <= _348;
        else
            _349 <= _346;
    end
    always @(posedge _84) begin
        if (_82)
            _352 <= _351;
        else
            _352 <= _349;
    end
    always @(posedge _84) begin
        if (_82)
            _355 <= _354;
        else
            _355 <= _352;
    end
    assign _356 = ~ _355;
    always @(posedge _84) begin
        if (_82)
            _304 <= _303;
        else
            _304 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _307 <= _306;
        else
            _307 <= _304;
    end
    always @(posedge _84) begin
        if (_82)
            _310 <= _309;
        else
            _310 <= _307;
    end
    always @(posedge _84) begin
        if (_82)
            _313 <= _312;
        else
            _313 <= _310;
    end
    always @(posedge _84) begin
        if (_82)
            _316 <= _315;
        else
            _316 <= _313;
    end
    always @(posedge _84) begin
        if (_82)
            _319 <= _318;
        else
            _319 <= _316;
    end
    always @(posedge _84) begin
        if (_82)
            _322 <= _321;
        else
            _322 <= _319;
    end
    always @(posedge _84) begin
        if (_82)
            _325 <= _324;
        else
            _325 <= _322;
    end
    always @(posedge _84) begin
        if (_82)
            _328 <= _327;
        else
            _328 <= _325;
    end
    assign _357 = _328 & _356;
    assign _358 = _129 & _357;
    assign write_enable_10 = _358 & PHASE_1;
    assign _363 = write_enable_10 | read_enable_8;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_4
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_363), .regcea(vdd), .wea(write_enable_10), .addra(address_10), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_1), .regceb(vdd), .web(write_enable_1), .addrb(address_1), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_370[131:131]), .sbiterrb(_370[130:130]), .doutb(_370[129:66]), .dbiterra(_370[65:65]), .sbiterra(_370[64:64]), .douta(_370[63:0]) );
    assign _371 = _370[63:0];
    assign _301 = ~ PHASE_1;
    assign _7 = _301;
    always @(posedge _84) begin
        if (_82)
            PHASE_1 <= _299;
        else
            if (_72)
                PHASE_1 <= _7;
    end
    assign _383 = PHASE_1 ? _382 : _371;
    assign address_11 = _568 ? _199 : _563;
    assign write_enable_11 = _561 & _568;
    assign address_12 = _568 ? _164 : _68;
    assign _570 = ~ _568;
    assign read_enable_9 = _556 & _570;
    assign _568 = ~ PHASE_4;
    assign write_enable_12 = _554 & _568;
    assign _572 = write_enable_12 | read_enable_9;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_5
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_572), .regcea(vdd), .wea(write_enable_12), .addra(address_12), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_11), .regceb(vdd), .web(write_enable_11), .addrb(address_11), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_577[131:131]), .sbiterrb(_577[130:130]), .doutb(_577[129:66]), .dbiterra(_577[65:65]), .sbiterra(_577[64:64]), .douta(_577[63:0]) );
    assign _578 = _577[63:0];
    assign address_13 = PHASE_4 ? _199 : _563;
    assign _561 = _129 & _524;
    assign write_enable_13 = _561 & PHASE_4;
    assign _486 = _478[129:66];
    assign _485 = _465[129:66];
    assign _487 = PHASE_2 ? _486 : _485;
    assign _483 = _423[129:66];
    assign _482 = _409[129:66];
    assign q1_0 = PHASE_3 ? _483 : _482;
    assign _488 = _390 ? _487 : q1_0;
    assign address_14 = _467 ? _461 : _460;
    assign _473 = ~ _467;
    assign read_enable_10 = _102 & _473;
    assign address_15 = _467 ? _60 : _443;
    assign _469 = ~ _467;
    assign read_enable_11 = _102 & _469;
    assign _467 = ~ PHASE_2;
    assign write_enable_15 = _426 & _467;
    assign _471 = write_enable_15 | read_enable_11;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_6
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_471), .regcea(vdd), .wea(write_enable_15), .addra(address_15), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_10), .regceb(vdd), .web(write_enable_14), .addrb(address_14), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_478[131:131]), .sbiterrb(_478[130:130]), .doutb(_478[129:66]), .dbiterra(_478[65:65]), .sbiterra(_478[64:64]), .douta(_478[63:0]) );
    assign _479 = _478[63:0];
    assign _459 = _172[11:11];
    assign _458 = _172[10:10];
    assign _457 = _172[9:9];
    assign _456 = _172[8:8];
    assign _455 = _172[7:7];
    assign _454 = _172[6:6];
    assign _453 = _172[5:5];
    assign _452 = _172[4:4];
    assign _451 = _172[3:3];
    assign _450 = _172[2:2];
    assign _449 = _172[1:1];
    assign _448 = _172[0:0];
    assign _460 = { _448, _449, _450, _451, _452, _453, _454, _455, _456, _457, _458, _459 };
    assign address_16 = PHASE_2 ? _461 : _460;
    assign _445 = ~ PHASE_2;
    assign read_enable_12 = _102 & _445;
    assign data_13 = wr_d6;
    assign _442 = _137[11:11];
    assign _441 = _137[10:10];
    assign _440 = _137[9:9];
    assign _439 = _137[8:8];
    assign _438 = _137[7:7];
    assign _437 = _137[6:6];
    assign _436 = _137[5:5];
    assign _435 = _137[4:4];
    assign _434 = _137[3:3];
    assign _433 = _137[2:2];
    assign _432 = _137[1:1];
    assign _431 = _137[0:0];
    assign _443 = { _431, _432, _433, _434, _435, _436, _437, _438, _439, _440, _441, _442 };
    assign address_17 = PHASE_2 ? _60 : _443;
    assign _428 = ~ PHASE_2;
    assign read_enable_13 = _102 & _428;
    assign _426 = _62[6:6];
    assign write_enable_17 = _426 & PHASE_2;
    assign _430 = write_enable_17 | read_enable_13;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_7
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_430), .regcea(vdd), .wea(write_enable_17), .addra(address_17), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_12), .regceb(vdd), .web(write_enable_16), .addrb(address_16), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_465[131:131]), .sbiterrb(_465[130:130]), .doutb(_465[129:66]), .dbiterra(_465[65:65]), .sbiterra(_465[64:64]), .douta(_465[63:0]) );
    assign _466 = _465[63:0];
    assign _387 = ~ PHASE_2;
    assign _11 = _387;
    always @(posedge _84) begin
        if (_82)
            PHASE_2 <= _385;
        else
            if (_72)
                PHASE_2 <= _11;
    end
    assign _480 = PHASE_2 ? _479 : _466;
    assign address_18 = _411 ? _199 : _172;
    assign _418 = ~ _411;
    assign read_enable_14 = _102 & _418;
    assign write_enable_18 = _402 & _411;
    assign _420 = write_enable_18 | read_enable_14;
    assign address_19 = _411 ? _164 : _137;
    assign _413 = ~ _411;
    assign read_enable_15 = _102 & _413;
    assign _411 = ~ PHASE_3;
    assign write_enable_19 = _395 & _411;
    assign _415 = write_enable_19 | read_enable_15;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_8
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_415), .regcea(vdd), .wea(write_enable_19), .addra(address_19), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_420), .regceb(vdd), .web(write_enable_18), .addrb(address_18), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_423[131:131]), .sbiterrb(_423[130:130]), .doutb(_423[129:66]), .dbiterra(_423[65:65]), .sbiterra(_423[64:64]), .douta(_423[63:0]) );
    assign _424 = _423[63:0];
    assign _491 = _490[127:64];
    assign data_15 = _491;
    assign address_20 = PHASE_3 ? _199 : _172;
    assign _404 = ~ PHASE_3;
    assign read_enable_16 = _102 & _404;
    assign _401 = ~ _130;
    assign _402 = _129 & _401;
    assign write_enable_20 = _402 & PHASE_3;
    assign _406 = write_enable_20 | read_enable_16;
    assign address_21 = PHASE_3 ? _164 : _137;
    assign _397 = ~ PHASE_3;
    assign read_enable_17 = _102 & _397;
    assign _394 = ~ _130;
    assign _395 = _129 & _394;
    assign write_enable_21 = _395 & PHASE_3;
    assign _399 = write_enable_21 | read_enable_17;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_9
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_399), .regcea(vdd), .wea(write_enable_21), .addra(address_21), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_406), .regceb(vdd), .web(write_enable_20), .addrb(address_20), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_409[131:131]), .sbiterrb(_409[130:130]), .doutb(_409[129:66]), .dbiterra(_409[65:65]), .sbiterra(_409[64:64]), .douta(_409[63:0]) );
    assign _410 = _409[63:0];
    assign _492 = ~ PHASE_3;
    assign _13 = _492;
    always @(posedge _84) begin
        if (_82)
            PHASE_3 <= _392;
        else
            if (_99)
                PHASE_3 <= _13;
    end
    assign q0_0 = PHASE_3 ? _424 : _410;
    always @(posedge _84) begin
        if (_82)
            _390 <= _389;
        else
            _390 <= _92;
    end
    assign _481 = _390 ? _480 : q0_0;
    dp_45
        dp_5
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_481), .d2(_488), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_490[191:128]), .q2(_490[127:64]), .q1(_490[63:0]) );
    assign _493 = _490[63:0];
    assign data_19 = _493;
    assign address_22 = PHASE_4 ? _164 : _68;
    assign _557 = ~ PHASE_4;
    assign _556 = _70[6:6];
    assign read_enable_18 = _556 & _557;
    always @(posedge _84) begin
        if (_82)
            _527 <= _526;
        else
            _527 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _530 <= _529;
        else
            _530 <= _527;
    end
    always @(posedge _84) begin
        if (_82)
            _533 <= _532;
        else
            _533 <= _530;
    end
    always @(posedge _84) begin
        if (_82)
            _536 <= _535;
        else
            _536 <= _533;
    end
    always @(posedge _84) begin
        if (_82)
            _539 <= _538;
        else
            _539 <= _536;
    end
    always @(posedge _84) begin
        if (_82)
            _542 <= _541;
        else
            _542 <= _539;
    end
    always @(posedge _84) begin
        if (_82)
            _545 <= _544;
        else
            _545 <= _542;
    end
    always @(posedge _84) begin
        if (_82)
            _548 <= _547;
        else
            _548 <= _545;
    end
    always @(posedge _84) begin
        if (_82)
            _551 <= _550;
        else
            _551 <= _548;
    end
    assign _552 = ~ _551;
    always @(posedge _84) begin
        if (_82)
            _500 <= _499;
        else
            _500 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _503 <= _502;
        else
            _503 <= _500;
    end
    always @(posedge _84) begin
        if (_82)
            _506 <= _505;
        else
            _506 <= _503;
    end
    always @(posedge _84) begin
        if (_82)
            _509 <= _508;
        else
            _509 <= _506;
    end
    always @(posedge _84) begin
        if (_82)
            _512 <= _511;
        else
            _512 <= _509;
    end
    always @(posedge _84) begin
        if (_82)
            _515 <= _514;
        else
            _515 <= _512;
    end
    always @(posedge _84) begin
        if (_82)
            _518 <= _517;
        else
            _518 <= _515;
    end
    always @(posedge _84) begin
        if (_82)
            _521 <= _520;
        else
            _521 <= _518;
    end
    always @(posedge _84) begin
        if (_82)
            _524 <= _523;
        else
            _524 <= _521;
    end
    assign _553 = _524 & _552;
    assign _554 = _129 & _553;
    assign write_enable_22 = _554 & PHASE_4;
    assign _559 = write_enable_22 | read_enable_18;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_10
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_559), .regcea(vdd), .wea(write_enable_22), .addra(address_22), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_13), .regceb(vdd), .web(write_enable_13), .addrb(address_13), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_566[131:131]), .sbiterrb(_566[130:130]), .doutb(_566[129:66]), .dbiterra(_566[65:65]), .sbiterra(_566[64:64]), .douta(_566[63:0]) );
    assign _567 = _566[63:0];
    assign _497 = ~ PHASE_4;
    assign _15 = _497;
    always @(posedge _84) begin
        if (_82)
            PHASE_4 <= _495;
        else
            if (_72)
                PHASE_4 <= _15;
    end
    assign _579 = PHASE_4 ? _578 : _567;
    assign address_23 = _764 ? _199 : _759;
    assign write_enable_23 = _757 & _764;
    assign address_24 = _764 ? _164 : _68;
    assign _766 = ~ _764;
    assign read_enable_19 = _752 & _766;
    assign _764 = ~ PHASE_7;
    assign write_enable_24 = _750 & _764;
    assign _768 = write_enable_24 | read_enable_19;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_11
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_768), .regcea(vdd), .wea(write_enable_24), .addra(address_24), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_23), .regceb(vdd), .web(write_enable_23), .addrb(address_23), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_773[131:131]), .sbiterrb(_773[130:130]), .doutb(_773[129:66]), .dbiterra(_773[65:65]), .sbiterra(_773[64:64]), .douta(_773[63:0]) );
    assign _774 = _773[63:0];
    assign address_25 = PHASE_7 ? _199 : _759;
    assign _757 = _129 & _720;
    assign write_enable_25 = _757 & PHASE_7;
    assign _682 = _674[129:66];
    assign _681 = _661[129:66];
    assign _683 = PHASE_5 ? _682 : _681;
    assign _679 = _619[129:66];
    assign _678 = _605[129:66];
    assign q1_1 = PHASE_6 ? _679 : _678;
    assign _684 = _586 ? _683 : q1_1;
    assign address_26 = _663 ? _657 : _656;
    assign _669 = ~ _663;
    assign read_enable_20 = _102 & _669;
    assign address_27 = _663 ? _60 : _639;
    assign _665 = ~ _663;
    assign read_enable_21 = _102 & _665;
    assign _663 = ~ PHASE_5;
    assign write_enable_27 = _622 & _663;
    assign _667 = write_enable_27 | read_enable_21;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_12
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_667), .regcea(vdd), .wea(write_enable_27), .addra(address_27), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_20), .regceb(vdd), .web(write_enable_26), .addrb(address_26), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_674[131:131]), .sbiterrb(_674[130:130]), .doutb(_674[129:66]), .dbiterra(_674[65:65]), .sbiterra(_674[64:64]), .douta(_674[63:0]) );
    assign _675 = _674[63:0];
    assign _655 = _172[11:11];
    assign _654 = _172[10:10];
    assign _653 = _172[9:9];
    assign _652 = _172[8:8];
    assign _651 = _172[7:7];
    assign _650 = _172[6:6];
    assign _649 = _172[5:5];
    assign _648 = _172[4:4];
    assign _647 = _172[3:3];
    assign _646 = _172[2:2];
    assign _645 = _172[1:1];
    assign _644 = _172[0:0];
    assign _656 = { _644, _645, _646, _647, _648, _649, _650, _651, _652, _653, _654, _655 };
    assign address_28 = PHASE_5 ? _657 : _656;
    assign _641 = ~ PHASE_5;
    assign read_enable_22 = _102 & _641;
    assign data_25 = wr_d5;
    assign _638 = _137[11:11];
    assign _637 = _137[10:10];
    assign _636 = _137[9:9];
    assign _635 = _137[8:8];
    assign _634 = _137[7:7];
    assign _633 = _137[6:6];
    assign _632 = _137[5:5];
    assign _631 = _137[4:4];
    assign _630 = _137[3:3];
    assign _629 = _137[2:2];
    assign _628 = _137[1:1];
    assign _627 = _137[0:0];
    assign _639 = { _627, _628, _629, _630, _631, _632, _633, _634, _635, _636, _637, _638 };
    assign address_29 = PHASE_5 ? _60 : _639;
    assign _624 = ~ PHASE_5;
    assign read_enable_23 = _102 & _624;
    assign _622 = _62[5:5];
    assign write_enable_29 = _622 & PHASE_5;
    assign _626 = write_enable_29 | read_enable_23;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_13
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_626), .regcea(vdd), .wea(write_enable_29), .addra(address_29), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_22), .regceb(vdd), .web(write_enable_28), .addrb(address_28), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_661[131:131]), .sbiterrb(_661[130:130]), .doutb(_661[129:66]), .dbiterra(_661[65:65]), .sbiterra(_661[64:64]), .douta(_661[63:0]) );
    assign _662 = _661[63:0];
    assign _583 = ~ PHASE_5;
    assign _19 = _583;
    always @(posedge _84) begin
        if (_82)
            PHASE_5 <= _581;
        else
            if (_72)
                PHASE_5 <= _19;
    end
    assign _676 = PHASE_5 ? _675 : _662;
    assign address_30 = _607 ? _199 : _172;
    assign _614 = ~ _607;
    assign read_enable_24 = _102 & _614;
    assign write_enable_30 = _598 & _607;
    assign _616 = write_enable_30 | read_enable_24;
    assign address_31 = _607 ? _164 : _137;
    assign _609 = ~ _607;
    assign read_enable_25 = _102 & _609;
    assign _607 = ~ PHASE_6;
    assign write_enable_31 = _591 & _607;
    assign _611 = write_enable_31 | read_enable_25;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_14
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_611), .regcea(vdd), .wea(write_enable_31), .addra(address_31), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_616), .regceb(vdd), .web(write_enable_30), .addrb(address_30), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_619[131:131]), .sbiterrb(_619[130:130]), .doutb(_619[129:66]), .dbiterra(_619[65:65]), .sbiterra(_619[64:64]), .douta(_619[63:0]) );
    assign _620 = _619[63:0];
    assign _687 = _686[127:64];
    assign data_27 = _687;
    assign address_32 = PHASE_6 ? _199 : _172;
    assign _600 = ~ PHASE_6;
    assign read_enable_26 = _102 & _600;
    assign _597 = ~ _130;
    assign _598 = _129 & _597;
    assign write_enable_32 = _598 & PHASE_6;
    assign _602 = write_enable_32 | read_enable_26;
    assign address_33 = PHASE_6 ? _164 : _137;
    assign _593 = ~ PHASE_6;
    assign read_enable_27 = _102 & _593;
    assign _590 = ~ _130;
    assign _591 = _129 & _590;
    assign write_enable_33 = _591 & PHASE_6;
    assign _595 = write_enable_33 | read_enable_27;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_15
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_595), .regcea(vdd), .wea(write_enable_33), .addra(address_33), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_602), .regceb(vdd), .web(write_enable_32), .addrb(address_32), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_605[131:131]), .sbiterrb(_605[130:130]), .doutb(_605[129:66]), .dbiterra(_605[65:65]), .sbiterra(_605[64:64]), .douta(_605[63:0]) );
    assign _606 = _605[63:0];
    assign _688 = ~ PHASE_6;
    assign _21 = _688;
    always @(posedge _84) begin
        if (_82)
            PHASE_6 <= _588;
        else
            if (_99)
                PHASE_6 <= _21;
    end
    assign q0_1 = PHASE_6 ? _620 : _606;
    always @(posedge _84) begin
        if (_82)
            _586 <= _585;
        else
            _586 <= _92;
    end
    assign _677 = _586 ? _676 : q0_1;
    dp_44
        dp_4
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_677), .d2(_684), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_686[191:128]), .q2(_686[127:64]), .q1(_686[63:0]) );
    assign _689 = _686[63:0];
    assign data_31 = _689;
    assign address_34 = PHASE_7 ? _164 : _68;
    assign _753 = ~ PHASE_7;
    assign _752 = _70[5:5];
    assign read_enable_28 = _752 & _753;
    always @(posedge _84) begin
        if (_82)
            _723 <= _722;
        else
            _723 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _726 <= _725;
        else
            _726 <= _723;
    end
    always @(posedge _84) begin
        if (_82)
            _729 <= _728;
        else
            _729 <= _726;
    end
    always @(posedge _84) begin
        if (_82)
            _732 <= _731;
        else
            _732 <= _729;
    end
    always @(posedge _84) begin
        if (_82)
            _735 <= _734;
        else
            _735 <= _732;
    end
    always @(posedge _84) begin
        if (_82)
            _738 <= _737;
        else
            _738 <= _735;
    end
    always @(posedge _84) begin
        if (_82)
            _741 <= _740;
        else
            _741 <= _738;
    end
    always @(posedge _84) begin
        if (_82)
            _744 <= _743;
        else
            _744 <= _741;
    end
    always @(posedge _84) begin
        if (_82)
            _747 <= _746;
        else
            _747 <= _744;
    end
    assign _748 = ~ _747;
    always @(posedge _84) begin
        if (_82)
            _696 <= _695;
        else
            _696 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _699 <= _698;
        else
            _699 <= _696;
    end
    always @(posedge _84) begin
        if (_82)
            _702 <= _701;
        else
            _702 <= _699;
    end
    always @(posedge _84) begin
        if (_82)
            _705 <= _704;
        else
            _705 <= _702;
    end
    always @(posedge _84) begin
        if (_82)
            _708 <= _707;
        else
            _708 <= _705;
    end
    always @(posedge _84) begin
        if (_82)
            _711 <= _710;
        else
            _711 <= _708;
    end
    always @(posedge _84) begin
        if (_82)
            _714 <= _713;
        else
            _714 <= _711;
    end
    always @(posedge _84) begin
        if (_82)
            _717 <= _716;
        else
            _717 <= _714;
    end
    always @(posedge _84) begin
        if (_82)
            _720 <= _719;
        else
            _720 <= _717;
    end
    assign _749 = _720 & _748;
    assign _750 = _129 & _749;
    assign write_enable_34 = _750 & PHASE_7;
    assign _755 = write_enable_34 | read_enable_28;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_16
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_755), .regcea(vdd), .wea(write_enable_34), .addra(address_34), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_25), .regceb(vdd), .web(write_enable_25), .addrb(address_25), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_762[131:131]), .sbiterrb(_762[130:130]), .doutb(_762[129:66]), .dbiterra(_762[65:65]), .sbiterra(_762[64:64]), .douta(_762[63:0]) );
    assign _763 = _762[63:0];
    assign _693 = ~ PHASE_7;
    assign _23 = _693;
    always @(posedge _84) begin
        if (_82)
            PHASE_7 <= _691;
        else
            if (_72)
                PHASE_7 <= _23;
    end
    assign _775 = PHASE_7 ? _774 : _763;
    assign address_35 = _960 ? _199 : _955;
    assign write_enable_35 = _953 & _960;
    assign address_36 = _960 ? _164 : _68;
    assign _962 = ~ _960;
    assign read_enable_29 = _948 & _962;
    assign _960 = ~ PHASE_10;
    assign write_enable_36 = _946 & _960;
    assign _964 = write_enable_36 | read_enable_29;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_17
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_964), .regcea(vdd), .wea(write_enable_36), .addra(address_36), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_35), .regceb(vdd), .web(write_enable_35), .addrb(address_35), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_969[131:131]), .sbiterrb(_969[130:130]), .doutb(_969[129:66]), .dbiterra(_969[65:65]), .sbiterra(_969[64:64]), .douta(_969[63:0]) );
    assign _970 = _969[63:0];
    assign address_37 = PHASE_10 ? _199 : _955;
    assign _953 = _129 & _916;
    assign write_enable_37 = _953 & PHASE_10;
    assign _878 = _870[129:66];
    assign _877 = _857[129:66];
    assign _879 = PHASE_8 ? _878 : _877;
    assign _875 = _815[129:66];
    assign _874 = _801[129:66];
    assign q1_2 = PHASE_9 ? _875 : _874;
    assign _880 = _782 ? _879 : q1_2;
    assign address_38 = _859 ? _853 : _852;
    assign _865 = ~ _859;
    assign read_enable_30 = _102 & _865;
    assign address_39 = _859 ? _60 : _835;
    assign _861 = ~ _859;
    assign read_enable_31 = _102 & _861;
    assign _859 = ~ PHASE_8;
    assign write_enable_39 = _818 & _859;
    assign _863 = write_enable_39 | read_enable_31;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_18
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_863), .regcea(vdd), .wea(write_enable_39), .addra(address_39), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_30), .regceb(vdd), .web(write_enable_38), .addrb(address_38), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_870[131:131]), .sbiterrb(_870[130:130]), .doutb(_870[129:66]), .dbiterra(_870[65:65]), .sbiterra(_870[64:64]), .douta(_870[63:0]) );
    assign _871 = _870[63:0];
    assign _851 = _172[11:11];
    assign _850 = _172[10:10];
    assign _849 = _172[9:9];
    assign _848 = _172[8:8];
    assign _847 = _172[7:7];
    assign _846 = _172[6:6];
    assign _845 = _172[5:5];
    assign _844 = _172[4:4];
    assign _843 = _172[3:3];
    assign _842 = _172[2:2];
    assign _841 = _172[1:1];
    assign _840 = _172[0:0];
    assign _852 = { _840, _841, _842, _843, _844, _845, _846, _847, _848, _849, _850, _851 };
    assign address_40 = PHASE_8 ? _853 : _852;
    assign _837 = ~ PHASE_8;
    assign read_enable_32 = _102 & _837;
    assign data_37 = wr_d4;
    assign _834 = _137[11:11];
    assign _833 = _137[10:10];
    assign _832 = _137[9:9];
    assign _831 = _137[8:8];
    assign _830 = _137[7:7];
    assign _829 = _137[6:6];
    assign _828 = _137[5:5];
    assign _827 = _137[4:4];
    assign _826 = _137[3:3];
    assign _825 = _137[2:2];
    assign _824 = _137[1:1];
    assign _823 = _137[0:0];
    assign _835 = { _823, _824, _825, _826, _827, _828, _829, _830, _831, _832, _833, _834 };
    assign address_41 = PHASE_8 ? _60 : _835;
    assign _820 = ~ PHASE_8;
    assign read_enable_33 = _102 & _820;
    assign _818 = _62[4:4];
    assign write_enable_41 = _818 & PHASE_8;
    assign _822 = write_enable_41 | read_enable_33;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_19
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_822), .regcea(vdd), .wea(write_enable_41), .addra(address_41), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_32), .regceb(vdd), .web(write_enable_40), .addrb(address_40), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_857[131:131]), .sbiterrb(_857[130:130]), .doutb(_857[129:66]), .dbiterra(_857[65:65]), .sbiterra(_857[64:64]), .douta(_857[63:0]) );
    assign _858 = _857[63:0];
    assign _779 = ~ PHASE_8;
    assign _27 = _779;
    always @(posedge _84) begin
        if (_82)
            PHASE_8 <= _777;
        else
            if (_72)
                PHASE_8 <= _27;
    end
    assign _872 = PHASE_8 ? _871 : _858;
    assign address_42 = _803 ? _199 : _172;
    assign _810 = ~ _803;
    assign read_enable_34 = _102 & _810;
    assign write_enable_42 = _794 & _803;
    assign _812 = write_enable_42 | read_enable_34;
    assign address_43 = _803 ? _164 : _137;
    assign _805 = ~ _803;
    assign read_enable_35 = _102 & _805;
    assign _803 = ~ PHASE_9;
    assign write_enable_43 = _787 & _803;
    assign _807 = write_enable_43 | read_enable_35;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_20
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_807), .regcea(vdd), .wea(write_enable_43), .addra(address_43), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_812), .regceb(vdd), .web(write_enable_42), .addrb(address_42), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_815[131:131]), .sbiterrb(_815[130:130]), .doutb(_815[129:66]), .dbiterra(_815[65:65]), .sbiterra(_815[64:64]), .douta(_815[63:0]) );
    assign _816 = _815[63:0];
    assign _883 = _882[127:64];
    assign data_39 = _883;
    assign address_44 = PHASE_9 ? _199 : _172;
    assign _796 = ~ PHASE_9;
    assign read_enable_36 = _102 & _796;
    assign _793 = ~ _130;
    assign _794 = _129 & _793;
    assign write_enable_44 = _794 & PHASE_9;
    assign _798 = write_enable_44 | read_enable_36;
    assign address_45 = PHASE_9 ? _164 : _137;
    assign _789 = ~ PHASE_9;
    assign read_enable_37 = _102 & _789;
    assign _786 = ~ _130;
    assign _787 = _129 & _786;
    assign write_enable_45 = _787 & PHASE_9;
    assign _791 = write_enable_45 | read_enable_37;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_21
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_791), .regcea(vdd), .wea(write_enable_45), .addra(address_45), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_798), .regceb(vdd), .web(write_enable_44), .addrb(address_44), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_801[131:131]), .sbiterrb(_801[130:130]), .doutb(_801[129:66]), .dbiterra(_801[65:65]), .sbiterra(_801[64:64]), .douta(_801[63:0]) );
    assign _802 = _801[63:0];
    assign _884 = ~ PHASE_9;
    assign _29 = _884;
    always @(posedge _84) begin
        if (_82)
            PHASE_9 <= _784;
        else
            if (_99)
                PHASE_9 <= _29;
    end
    assign q0_2 = PHASE_9 ? _816 : _802;
    always @(posedge _84) begin
        if (_82)
            _782 <= _781;
        else
            _782 <= _92;
    end
    assign _873 = _782 ? _872 : q0_2;
    dp_43
        dp_3
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_873), .d2(_880), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_882[191:128]), .q2(_882[127:64]), .q1(_882[63:0]) );
    assign _885 = _882[63:0];
    assign data_43 = _885;
    assign address_46 = PHASE_10 ? _164 : _68;
    assign _949 = ~ PHASE_10;
    assign _948 = _70[4:4];
    assign read_enable_38 = _948 & _949;
    always @(posedge _84) begin
        if (_82)
            _919 <= _918;
        else
            _919 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _922 <= _921;
        else
            _922 <= _919;
    end
    always @(posedge _84) begin
        if (_82)
            _925 <= _924;
        else
            _925 <= _922;
    end
    always @(posedge _84) begin
        if (_82)
            _928 <= _927;
        else
            _928 <= _925;
    end
    always @(posedge _84) begin
        if (_82)
            _931 <= _930;
        else
            _931 <= _928;
    end
    always @(posedge _84) begin
        if (_82)
            _934 <= _933;
        else
            _934 <= _931;
    end
    always @(posedge _84) begin
        if (_82)
            _937 <= _936;
        else
            _937 <= _934;
    end
    always @(posedge _84) begin
        if (_82)
            _940 <= _939;
        else
            _940 <= _937;
    end
    always @(posedge _84) begin
        if (_82)
            _943 <= _942;
        else
            _943 <= _940;
    end
    assign _944 = ~ _943;
    always @(posedge _84) begin
        if (_82)
            _892 <= _891;
        else
            _892 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _895 <= _894;
        else
            _895 <= _892;
    end
    always @(posedge _84) begin
        if (_82)
            _898 <= _897;
        else
            _898 <= _895;
    end
    always @(posedge _84) begin
        if (_82)
            _901 <= _900;
        else
            _901 <= _898;
    end
    always @(posedge _84) begin
        if (_82)
            _904 <= _903;
        else
            _904 <= _901;
    end
    always @(posedge _84) begin
        if (_82)
            _907 <= _906;
        else
            _907 <= _904;
    end
    always @(posedge _84) begin
        if (_82)
            _910 <= _909;
        else
            _910 <= _907;
    end
    always @(posedge _84) begin
        if (_82)
            _913 <= _912;
        else
            _913 <= _910;
    end
    always @(posedge _84) begin
        if (_82)
            _916 <= _915;
        else
            _916 <= _913;
    end
    assign _945 = _916 & _944;
    assign _946 = _129 & _945;
    assign write_enable_46 = _946 & PHASE_10;
    assign _951 = write_enable_46 | read_enable_38;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_22
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_951), .regcea(vdd), .wea(write_enable_46), .addra(address_46), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_37), .regceb(vdd), .web(write_enable_37), .addrb(address_37), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_958[131:131]), .sbiterrb(_958[130:130]), .doutb(_958[129:66]), .dbiterra(_958[65:65]), .sbiterra(_958[64:64]), .douta(_958[63:0]) );
    assign _959 = _958[63:0];
    assign _889 = ~ PHASE_10;
    assign _31 = _889;
    always @(posedge _84) begin
        if (_82)
            PHASE_10 <= _887;
        else
            if (_72)
                PHASE_10 <= _31;
    end
    assign _971 = PHASE_10 ? _970 : _959;
    assign address_47 = _1156 ? _199 : _1151;
    assign write_enable_47 = _1149 & _1156;
    assign address_48 = _1156 ? _164 : _68;
    assign _1158 = ~ _1156;
    assign read_enable_39 = _1144 & _1158;
    assign _1156 = ~ PHASE_13;
    assign write_enable_48 = _1142 & _1156;
    assign _1160 = write_enable_48 | read_enable_39;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_23
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1160), .regcea(vdd), .wea(write_enable_48), .addra(address_48), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_47), .regceb(vdd), .web(write_enable_47), .addrb(address_47), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1165[131:131]), .sbiterrb(_1165[130:130]), .doutb(_1165[129:66]), .dbiterra(_1165[65:65]), .sbiterra(_1165[64:64]), .douta(_1165[63:0]) );
    assign _1166 = _1165[63:0];
    assign address_49 = PHASE_13 ? _199 : _1151;
    assign _1149 = _129 & _1112;
    assign write_enable_49 = _1149 & PHASE_13;
    assign _1074 = _1066[129:66];
    assign _1073 = _1053[129:66];
    assign _1075 = PHASE_11 ? _1074 : _1073;
    assign _1071 = _1011[129:66];
    assign _1070 = _997[129:66];
    assign q1_3 = PHASE_12 ? _1071 : _1070;
    assign _1076 = _978 ? _1075 : q1_3;
    assign address_50 = _1055 ? _1049 : _1048;
    assign _1061 = ~ _1055;
    assign read_enable_40 = _102 & _1061;
    assign address_51 = _1055 ? _60 : _1031;
    assign _1057 = ~ _1055;
    assign read_enable_41 = _102 & _1057;
    assign _1055 = ~ PHASE_11;
    assign write_enable_51 = _1014 & _1055;
    assign _1059 = write_enable_51 | read_enable_41;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_24
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1059), .regcea(vdd), .wea(write_enable_51), .addra(address_51), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_40), .regceb(vdd), .web(write_enable_50), .addrb(address_50), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1066[131:131]), .sbiterrb(_1066[130:130]), .doutb(_1066[129:66]), .dbiterra(_1066[65:65]), .sbiterra(_1066[64:64]), .douta(_1066[63:0]) );
    assign _1067 = _1066[63:0];
    assign _1047 = _172[11:11];
    assign _1046 = _172[10:10];
    assign _1045 = _172[9:9];
    assign _1044 = _172[8:8];
    assign _1043 = _172[7:7];
    assign _1042 = _172[6:6];
    assign _1041 = _172[5:5];
    assign _1040 = _172[4:4];
    assign _1039 = _172[3:3];
    assign _1038 = _172[2:2];
    assign _1037 = _172[1:1];
    assign _1036 = _172[0:0];
    assign _1048 = { _1036, _1037, _1038, _1039, _1040, _1041, _1042, _1043, _1044, _1045, _1046, _1047 };
    assign address_52 = PHASE_11 ? _1049 : _1048;
    assign _1033 = ~ PHASE_11;
    assign read_enable_42 = _102 & _1033;
    assign data_49 = wr_d3;
    assign _1030 = _137[11:11];
    assign _1029 = _137[10:10];
    assign _1028 = _137[9:9];
    assign _1027 = _137[8:8];
    assign _1026 = _137[7:7];
    assign _1025 = _137[6:6];
    assign _1024 = _137[5:5];
    assign _1023 = _137[4:4];
    assign _1022 = _137[3:3];
    assign _1021 = _137[2:2];
    assign _1020 = _137[1:1];
    assign _1019 = _137[0:0];
    assign _1031 = { _1019, _1020, _1021, _1022, _1023, _1024, _1025, _1026, _1027, _1028, _1029, _1030 };
    assign address_53 = PHASE_11 ? _60 : _1031;
    assign _1016 = ~ PHASE_11;
    assign read_enable_43 = _102 & _1016;
    assign _1014 = _62[3:3];
    assign write_enable_53 = _1014 & PHASE_11;
    assign _1018 = write_enable_53 | read_enable_43;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_25
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1018), .regcea(vdd), .wea(write_enable_53), .addra(address_53), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_42), .regceb(vdd), .web(write_enable_52), .addrb(address_52), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1053[131:131]), .sbiterrb(_1053[130:130]), .doutb(_1053[129:66]), .dbiterra(_1053[65:65]), .sbiterra(_1053[64:64]), .douta(_1053[63:0]) );
    assign _1054 = _1053[63:0];
    assign _975 = ~ PHASE_11;
    assign _35 = _975;
    always @(posedge _84) begin
        if (_82)
            PHASE_11 <= _973;
        else
            if (_72)
                PHASE_11 <= _35;
    end
    assign _1068 = PHASE_11 ? _1067 : _1054;
    assign address_54 = _999 ? _199 : _172;
    assign _1006 = ~ _999;
    assign read_enable_44 = _102 & _1006;
    assign write_enable_54 = _990 & _999;
    assign _1008 = write_enable_54 | read_enable_44;
    assign address_55 = _999 ? _164 : _137;
    assign _1001 = ~ _999;
    assign read_enable_45 = _102 & _1001;
    assign _999 = ~ PHASE_12;
    assign write_enable_55 = _983 & _999;
    assign _1003 = write_enable_55 | read_enable_45;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_26
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1003), .regcea(vdd), .wea(write_enable_55), .addra(address_55), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1008), .regceb(vdd), .web(write_enable_54), .addrb(address_54), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1011[131:131]), .sbiterrb(_1011[130:130]), .doutb(_1011[129:66]), .dbiterra(_1011[65:65]), .sbiterra(_1011[64:64]), .douta(_1011[63:0]) );
    assign _1012 = _1011[63:0];
    assign _1079 = _1078[127:64];
    assign data_51 = _1079;
    assign address_56 = PHASE_12 ? _199 : _172;
    assign _992 = ~ PHASE_12;
    assign read_enable_46 = _102 & _992;
    assign _989 = ~ _130;
    assign _990 = _129 & _989;
    assign write_enable_56 = _990 & PHASE_12;
    assign _994 = write_enable_56 | read_enable_46;
    assign address_57 = PHASE_12 ? _164 : _137;
    assign _985 = ~ PHASE_12;
    assign read_enable_47 = _102 & _985;
    assign _982 = ~ _130;
    assign _983 = _129 & _982;
    assign write_enable_57 = _983 & PHASE_12;
    assign _987 = write_enable_57 | read_enable_47;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_27
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_987), .regcea(vdd), .wea(write_enable_57), .addra(address_57), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_994), .regceb(vdd), .web(write_enable_56), .addrb(address_56), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_997[131:131]), .sbiterrb(_997[130:130]), .doutb(_997[129:66]), .dbiterra(_997[65:65]), .sbiterra(_997[64:64]), .douta(_997[63:0]) );
    assign _998 = _997[63:0];
    assign _1080 = ~ PHASE_12;
    assign _37 = _1080;
    always @(posedge _84) begin
        if (_82)
            PHASE_12 <= _980;
        else
            if (_99)
                PHASE_12 <= _37;
    end
    assign q0_3 = PHASE_12 ? _1012 : _998;
    always @(posedge _84) begin
        if (_82)
            _978 <= _977;
        else
            _978 <= _92;
    end
    assign _1069 = _978 ? _1068 : q0_3;
    dp_42
        dp_2
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1069), .d2(_1076), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1078[191:128]), .q2(_1078[127:64]), .q1(_1078[63:0]) );
    assign _1081 = _1078[63:0];
    assign data_55 = _1081;
    assign address_58 = PHASE_13 ? _164 : _68;
    assign _1145 = ~ PHASE_13;
    assign _1144 = _70[3:3];
    assign read_enable_48 = _1144 & _1145;
    always @(posedge _84) begin
        if (_82)
            _1115 <= _1114;
        else
            _1115 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1118 <= _1117;
        else
            _1118 <= _1115;
    end
    always @(posedge _84) begin
        if (_82)
            _1121 <= _1120;
        else
            _1121 <= _1118;
    end
    always @(posedge _84) begin
        if (_82)
            _1124 <= _1123;
        else
            _1124 <= _1121;
    end
    always @(posedge _84) begin
        if (_82)
            _1127 <= _1126;
        else
            _1127 <= _1124;
    end
    always @(posedge _84) begin
        if (_82)
            _1130 <= _1129;
        else
            _1130 <= _1127;
    end
    always @(posedge _84) begin
        if (_82)
            _1133 <= _1132;
        else
            _1133 <= _1130;
    end
    always @(posedge _84) begin
        if (_82)
            _1136 <= _1135;
        else
            _1136 <= _1133;
    end
    always @(posedge _84) begin
        if (_82)
            _1139 <= _1138;
        else
            _1139 <= _1136;
    end
    assign _1140 = ~ _1139;
    always @(posedge _84) begin
        if (_82)
            _1088 <= _1087;
        else
            _1088 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1091 <= _1090;
        else
            _1091 <= _1088;
    end
    always @(posedge _84) begin
        if (_82)
            _1094 <= _1093;
        else
            _1094 <= _1091;
    end
    always @(posedge _84) begin
        if (_82)
            _1097 <= _1096;
        else
            _1097 <= _1094;
    end
    always @(posedge _84) begin
        if (_82)
            _1100 <= _1099;
        else
            _1100 <= _1097;
    end
    always @(posedge _84) begin
        if (_82)
            _1103 <= _1102;
        else
            _1103 <= _1100;
    end
    always @(posedge _84) begin
        if (_82)
            _1106 <= _1105;
        else
            _1106 <= _1103;
    end
    always @(posedge _84) begin
        if (_82)
            _1109 <= _1108;
        else
            _1109 <= _1106;
    end
    always @(posedge _84) begin
        if (_82)
            _1112 <= _1111;
        else
            _1112 <= _1109;
    end
    assign _1141 = _1112 & _1140;
    assign _1142 = _129 & _1141;
    assign write_enable_58 = _1142 & PHASE_13;
    assign _1147 = write_enable_58 | read_enable_48;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_28
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1147), .regcea(vdd), .wea(write_enable_58), .addra(address_58), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_49), .regceb(vdd), .web(write_enable_49), .addrb(address_49), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1154[131:131]), .sbiterrb(_1154[130:130]), .doutb(_1154[129:66]), .dbiterra(_1154[65:65]), .sbiterra(_1154[64:64]), .douta(_1154[63:0]) );
    assign _1155 = _1154[63:0];
    assign _1085 = ~ PHASE_13;
    assign _39 = _1085;
    always @(posedge _84) begin
        if (_82)
            PHASE_13 <= _1083;
        else
            if (_72)
                PHASE_13 <= _39;
    end
    assign _1167 = PHASE_13 ? _1166 : _1155;
    assign address_59 = _1352 ? _199 : _1347;
    assign write_enable_59 = _1345 & _1352;
    assign address_60 = _1352 ? _164 : _68;
    assign _1354 = ~ _1352;
    assign read_enable_49 = _1340 & _1354;
    assign _1352 = ~ PHASE_16;
    assign write_enable_60 = _1338 & _1352;
    assign _1356 = write_enable_60 | read_enable_49;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_29
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1356), .regcea(vdd), .wea(write_enable_60), .addra(address_60), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_59), .regceb(vdd), .web(write_enable_59), .addrb(address_59), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1361[131:131]), .sbiterrb(_1361[130:130]), .doutb(_1361[129:66]), .dbiterra(_1361[65:65]), .sbiterra(_1361[64:64]), .douta(_1361[63:0]) );
    assign _1362 = _1361[63:0];
    assign address_61 = PHASE_16 ? _199 : _1347;
    assign _1345 = _129 & _1308;
    assign write_enable_61 = _1345 & PHASE_16;
    assign _1270 = _1262[129:66];
    assign _1269 = _1249[129:66];
    assign _1271 = PHASE_14 ? _1270 : _1269;
    assign _1267 = _1207[129:66];
    assign _1266 = _1193[129:66];
    assign q1_4 = PHASE_15 ? _1267 : _1266;
    assign _1272 = _1174 ? _1271 : q1_4;
    assign address_62 = _1251 ? _1245 : _1244;
    assign _1257 = ~ _1251;
    assign read_enable_50 = _102 & _1257;
    assign address_63 = _1251 ? _60 : _1227;
    assign _1253 = ~ _1251;
    assign read_enable_51 = _102 & _1253;
    assign _1251 = ~ PHASE_14;
    assign write_enable_63 = _1210 & _1251;
    assign _1255 = write_enable_63 | read_enable_51;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_30
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1255), .regcea(vdd), .wea(write_enable_63), .addra(address_63), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_50), .regceb(vdd), .web(write_enable_62), .addrb(address_62), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1262[131:131]), .sbiterrb(_1262[130:130]), .doutb(_1262[129:66]), .dbiterra(_1262[65:65]), .sbiterra(_1262[64:64]), .douta(_1262[63:0]) );
    assign _1263 = _1262[63:0];
    assign _1243 = _172[11:11];
    assign _1242 = _172[10:10];
    assign _1241 = _172[9:9];
    assign _1240 = _172[8:8];
    assign _1239 = _172[7:7];
    assign _1238 = _172[6:6];
    assign _1237 = _172[5:5];
    assign _1236 = _172[4:4];
    assign _1235 = _172[3:3];
    assign _1234 = _172[2:2];
    assign _1233 = _172[1:1];
    assign _1232 = _172[0:0];
    assign _1244 = { _1232, _1233, _1234, _1235, _1236, _1237, _1238, _1239, _1240, _1241, _1242, _1243 };
    assign address_64 = PHASE_14 ? _1245 : _1244;
    assign _1229 = ~ PHASE_14;
    assign read_enable_52 = _102 & _1229;
    assign data_61 = wr_d2;
    assign _1226 = _137[11:11];
    assign _1225 = _137[10:10];
    assign _1224 = _137[9:9];
    assign _1223 = _137[8:8];
    assign _1222 = _137[7:7];
    assign _1221 = _137[6:6];
    assign _1220 = _137[5:5];
    assign _1219 = _137[4:4];
    assign _1218 = _137[3:3];
    assign _1217 = _137[2:2];
    assign _1216 = _137[1:1];
    assign _1215 = _137[0:0];
    assign _1227 = { _1215, _1216, _1217, _1218, _1219, _1220, _1221, _1222, _1223, _1224, _1225, _1226 };
    assign address_65 = PHASE_14 ? _60 : _1227;
    assign _1212 = ~ PHASE_14;
    assign read_enable_53 = _102 & _1212;
    assign _1210 = _62[2:2];
    assign write_enable_65 = _1210 & PHASE_14;
    assign _1214 = write_enable_65 | read_enable_53;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_31
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1214), .regcea(vdd), .wea(write_enable_65), .addra(address_65), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_52), .regceb(vdd), .web(write_enable_64), .addrb(address_64), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1249[131:131]), .sbiterrb(_1249[130:130]), .doutb(_1249[129:66]), .dbiterra(_1249[65:65]), .sbiterra(_1249[64:64]), .douta(_1249[63:0]) );
    assign _1250 = _1249[63:0];
    assign _1171 = ~ PHASE_14;
    assign _43 = _1171;
    always @(posedge _84) begin
        if (_82)
            PHASE_14 <= _1169;
        else
            if (_72)
                PHASE_14 <= _43;
    end
    assign _1264 = PHASE_14 ? _1263 : _1250;
    assign address_66 = _1195 ? _199 : _172;
    assign _1202 = ~ _1195;
    assign read_enable_54 = _102 & _1202;
    assign write_enable_66 = _1186 & _1195;
    assign _1204 = write_enable_66 | read_enable_54;
    assign address_67 = _1195 ? _164 : _137;
    assign _1197 = ~ _1195;
    assign read_enable_55 = _102 & _1197;
    assign _1195 = ~ PHASE_15;
    assign write_enable_67 = _1179 & _1195;
    assign _1199 = write_enable_67 | read_enable_55;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_32
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1199), .regcea(vdd), .wea(write_enable_67), .addra(address_67), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1204), .regceb(vdd), .web(write_enable_66), .addrb(address_66), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1207[131:131]), .sbiterrb(_1207[130:130]), .doutb(_1207[129:66]), .dbiterra(_1207[65:65]), .sbiterra(_1207[64:64]), .douta(_1207[63:0]) );
    assign _1208 = _1207[63:0];
    assign _1275 = _1274[127:64];
    assign data_63 = _1275;
    assign address_68 = PHASE_15 ? _199 : _172;
    assign _1188 = ~ PHASE_15;
    assign read_enable_56 = _102 & _1188;
    assign _1185 = ~ _130;
    assign _1186 = _129 & _1185;
    assign write_enable_68 = _1186 & PHASE_15;
    assign _1190 = write_enable_68 | read_enable_56;
    assign address_69 = PHASE_15 ? _164 : _137;
    assign _1181 = ~ PHASE_15;
    assign read_enable_57 = _102 & _1181;
    assign _1178 = ~ _130;
    assign _1179 = _129 & _1178;
    assign write_enable_69 = _1179 & PHASE_15;
    assign _1183 = write_enable_69 | read_enable_57;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_33
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1183), .regcea(vdd), .wea(write_enable_69), .addra(address_69), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1190), .regceb(vdd), .web(write_enable_68), .addrb(address_68), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1193[131:131]), .sbiterrb(_1193[130:130]), .doutb(_1193[129:66]), .dbiterra(_1193[65:65]), .sbiterra(_1193[64:64]), .douta(_1193[63:0]) );
    assign _1194 = _1193[63:0];
    assign _1276 = ~ PHASE_15;
    assign _45 = _1276;
    always @(posedge _84) begin
        if (_82)
            PHASE_15 <= _1176;
        else
            if (_99)
                PHASE_15 <= _45;
    end
    assign q0_4 = PHASE_15 ? _1208 : _1194;
    always @(posedge _84) begin
        if (_82)
            _1174 <= _1173;
        else
            _1174 <= _92;
    end
    assign _1265 = _1174 ? _1264 : q0_4;
    dp_41
        dp_1
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1265), .d2(_1272), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1274[191:128]), .q2(_1274[127:64]), .q1(_1274[63:0]) );
    assign _1277 = _1274[63:0];
    assign data_67 = _1277;
    assign address_70 = PHASE_16 ? _164 : _68;
    assign _1341 = ~ PHASE_16;
    assign _1340 = _70[2:2];
    assign read_enable_58 = _1340 & _1341;
    always @(posedge _84) begin
        if (_82)
            _1311 <= _1310;
        else
            _1311 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1314 <= _1313;
        else
            _1314 <= _1311;
    end
    always @(posedge _84) begin
        if (_82)
            _1317 <= _1316;
        else
            _1317 <= _1314;
    end
    always @(posedge _84) begin
        if (_82)
            _1320 <= _1319;
        else
            _1320 <= _1317;
    end
    always @(posedge _84) begin
        if (_82)
            _1323 <= _1322;
        else
            _1323 <= _1320;
    end
    always @(posedge _84) begin
        if (_82)
            _1326 <= _1325;
        else
            _1326 <= _1323;
    end
    always @(posedge _84) begin
        if (_82)
            _1329 <= _1328;
        else
            _1329 <= _1326;
    end
    always @(posedge _84) begin
        if (_82)
            _1332 <= _1331;
        else
            _1332 <= _1329;
    end
    always @(posedge _84) begin
        if (_82)
            _1335 <= _1334;
        else
            _1335 <= _1332;
    end
    assign _1336 = ~ _1335;
    always @(posedge _84) begin
        if (_82)
            _1284 <= _1283;
        else
            _1284 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1287 <= _1286;
        else
            _1287 <= _1284;
    end
    always @(posedge _84) begin
        if (_82)
            _1290 <= _1289;
        else
            _1290 <= _1287;
    end
    always @(posedge _84) begin
        if (_82)
            _1293 <= _1292;
        else
            _1293 <= _1290;
    end
    always @(posedge _84) begin
        if (_82)
            _1296 <= _1295;
        else
            _1296 <= _1293;
    end
    always @(posedge _84) begin
        if (_82)
            _1299 <= _1298;
        else
            _1299 <= _1296;
    end
    always @(posedge _84) begin
        if (_82)
            _1302 <= _1301;
        else
            _1302 <= _1299;
    end
    always @(posedge _84) begin
        if (_82)
            _1305 <= _1304;
        else
            _1305 <= _1302;
    end
    always @(posedge _84) begin
        if (_82)
            _1308 <= _1307;
        else
            _1308 <= _1305;
    end
    assign _1337 = _1308 & _1336;
    assign _1338 = _129 & _1337;
    assign write_enable_70 = _1338 & PHASE_16;
    assign _1343 = write_enable_70 | read_enable_58;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_34
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1343), .regcea(vdd), .wea(write_enable_70), .addra(address_70), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_61), .regceb(vdd), .web(write_enable_61), .addrb(address_61), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1350[131:131]), .sbiterrb(_1350[130:130]), .doutb(_1350[129:66]), .dbiterra(_1350[65:65]), .sbiterra(_1350[64:64]), .douta(_1350[63:0]) );
    assign _1351 = _1350[63:0];
    assign _1281 = ~ PHASE_16;
    assign _47 = _1281;
    always @(posedge _84) begin
        if (_82)
            PHASE_16 <= _1279;
        else
            if (_72)
                PHASE_16 <= _47;
    end
    assign _1363 = PHASE_16 ? _1362 : _1351;
    assign address_71 = _1548 ? _199 : _1543;
    assign write_enable_71 = _1541 & _1548;
    assign address_72 = _1548 ? _164 : _68;
    assign _1550 = ~ _1548;
    assign read_enable_59 = _1536 & _1550;
    assign _1548 = ~ PHASE_19;
    assign write_enable_72 = _1534 & _1548;
    assign _1552 = write_enable_72 | read_enable_59;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_35
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1552), .regcea(vdd), .wea(write_enable_72), .addra(address_72), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_71), .regceb(vdd), .web(write_enable_71), .addrb(address_71), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1557[131:131]), .sbiterrb(_1557[130:130]), .doutb(_1557[129:66]), .dbiterra(_1557[65:65]), .sbiterra(_1557[64:64]), .douta(_1557[63:0]) );
    assign _1558 = _1557[63:0];
    assign address_73 = PHASE_19 ? _199 : _1543;
    assign _1541 = _129 & _1504;
    assign write_enable_73 = _1541 & PHASE_19;
    assign _1466 = _1458[129:66];
    assign _1465 = _1445[129:66];
    assign _1467 = PHASE_17 ? _1466 : _1465;
    assign _1463 = _1403[129:66];
    assign _1462 = _1389[129:66];
    assign q1_5 = PHASE_18 ? _1463 : _1462;
    assign _1468 = _1370 ? _1467 : q1_5;
    assign address_74 = _1447 ? _1441 : _1440;
    assign _1453 = ~ _1447;
    assign read_enable_60 = _102 & _1453;
    assign address_75 = _1447 ? _60 : _1423;
    assign _1449 = ~ _1447;
    assign read_enable_61 = _102 & _1449;
    assign _1447 = ~ PHASE_17;
    assign write_enable_75 = _1406 & _1447;
    assign _1451 = write_enable_75 | read_enable_61;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_36
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1451), .regcea(vdd), .wea(write_enable_75), .addra(address_75), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_60), .regceb(vdd), .web(write_enable_74), .addrb(address_74), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1458[131:131]), .sbiterrb(_1458[130:130]), .doutb(_1458[129:66]), .dbiterra(_1458[65:65]), .sbiterra(_1458[64:64]), .douta(_1458[63:0]) );
    assign _1459 = _1458[63:0];
    assign _1439 = _172[11:11];
    assign _1438 = _172[10:10];
    assign _1437 = _172[9:9];
    assign _1436 = _172[8:8];
    assign _1435 = _172[7:7];
    assign _1434 = _172[6:6];
    assign _1433 = _172[5:5];
    assign _1432 = _172[4:4];
    assign _1431 = _172[3:3];
    assign _1430 = _172[2:2];
    assign _1429 = _172[1:1];
    assign _1428 = _172[0:0];
    assign _1440 = { _1428, _1429, _1430, _1431, _1432, _1433, _1434, _1435, _1436, _1437, _1438, _1439 };
    assign address_76 = PHASE_17 ? _1441 : _1440;
    assign _1425 = ~ PHASE_17;
    assign read_enable_62 = _102 & _1425;
    assign data_73 = wr_d1;
    assign _1422 = _137[11:11];
    assign _1421 = _137[10:10];
    assign _1420 = _137[9:9];
    assign _1419 = _137[8:8];
    assign _1418 = _137[7:7];
    assign _1417 = _137[6:6];
    assign _1416 = _137[5:5];
    assign _1415 = _137[4:4];
    assign _1414 = _137[3:3];
    assign _1413 = _137[2:2];
    assign _1412 = _137[1:1];
    assign _1411 = _137[0:0];
    assign _1423 = { _1411, _1412, _1413, _1414, _1415, _1416, _1417, _1418, _1419, _1420, _1421, _1422 };
    assign address_77 = PHASE_17 ? _60 : _1423;
    assign _1408 = ~ PHASE_17;
    assign read_enable_63 = _102 & _1408;
    assign _1406 = _62[1:1];
    assign write_enable_77 = _1406 & PHASE_17;
    assign _1410 = write_enable_77 | read_enable_63;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_37
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1410), .regcea(vdd), .wea(write_enable_77), .addra(address_77), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_62), .regceb(vdd), .web(write_enable_76), .addrb(address_76), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1445[131:131]), .sbiterrb(_1445[130:130]), .doutb(_1445[129:66]), .dbiterra(_1445[65:65]), .sbiterra(_1445[64:64]), .douta(_1445[63:0]) );
    assign _1446 = _1445[63:0];
    assign _1367 = ~ PHASE_17;
    assign _51 = _1367;
    always @(posedge _84) begin
        if (_82)
            PHASE_17 <= _1365;
        else
            if (_72)
                PHASE_17 <= _51;
    end
    assign _1460 = PHASE_17 ? _1459 : _1446;
    assign address_78 = _1391 ? _199 : _172;
    assign _1398 = ~ _1391;
    assign read_enable_64 = _102 & _1398;
    assign write_enable_78 = _1382 & _1391;
    assign _1400 = write_enable_78 | read_enable_64;
    assign address_79 = _1391 ? _164 : _137;
    assign _1393 = ~ _1391;
    assign read_enable_65 = _102 & _1393;
    assign _1391 = ~ PHASE_18;
    assign write_enable_79 = _1375 & _1391;
    assign _1395 = write_enable_79 | read_enable_65;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_38
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1395), .regcea(vdd), .wea(write_enable_79), .addra(address_79), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1400), .regceb(vdd), .web(write_enable_78), .addrb(address_78), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1403[131:131]), .sbiterrb(_1403[130:130]), .doutb(_1403[129:66]), .dbiterra(_1403[65:65]), .sbiterra(_1403[64:64]), .douta(_1403[63:0]) );
    assign _1404 = _1403[63:0];
    assign _1471 = _1470[127:64];
    assign data_75 = _1471;
    assign address_80 = PHASE_18 ? _199 : _172;
    assign _1384 = ~ PHASE_18;
    assign read_enable_66 = _102 & _1384;
    assign _1381 = ~ _130;
    assign _1382 = _129 & _1381;
    assign write_enable_80 = _1382 & PHASE_18;
    assign _1386 = write_enable_80 | read_enable_66;
    assign address_81 = PHASE_18 ? _164 : _137;
    assign _1377 = ~ PHASE_18;
    assign read_enable_67 = _102 & _1377;
    assign _1374 = ~ _130;
    assign _1375 = _129 & _1374;
    assign write_enable_81 = _1375 & PHASE_18;
    assign _1379 = write_enable_81 | read_enable_67;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_39
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1379), .regcea(vdd), .wea(write_enable_81), .addra(address_81), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1386), .regceb(vdd), .web(write_enable_80), .addrb(address_80), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1389[131:131]), .sbiterrb(_1389[130:130]), .doutb(_1389[129:66]), .dbiterra(_1389[65:65]), .sbiterra(_1389[64:64]), .douta(_1389[63:0]) );
    assign _1390 = _1389[63:0];
    assign _1472 = ~ PHASE_18;
    assign _53 = _1472;
    always @(posedge _84) begin
        if (_82)
            PHASE_18 <= _1372;
        else
            if (_99)
                PHASE_18 <= _53;
    end
    assign q0_5 = PHASE_18 ? _1404 : _1390;
    always @(posedge _84) begin
        if (_82)
            _1370 <= _1369;
        else
            _1370 <= _92;
    end
    assign _1461 = _1370 ? _1460 : q0_5;
    dp_40
        dp_0
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1461), .d2(_1468), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1470[191:128]), .q2(_1470[127:64]), .q1(_1470[63:0]) );
    assign _1473 = _1470[63:0];
    assign data_79 = _1473;
    assign address_82 = PHASE_19 ? _164 : _68;
    assign _1537 = ~ PHASE_19;
    assign _1536 = _70[1:1];
    assign read_enable_68 = _1536 & _1537;
    always @(posedge _84) begin
        if (_82)
            _1507 <= _1506;
        else
            _1507 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1510 <= _1509;
        else
            _1510 <= _1507;
    end
    always @(posedge _84) begin
        if (_82)
            _1513 <= _1512;
        else
            _1513 <= _1510;
    end
    always @(posedge _84) begin
        if (_82)
            _1516 <= _1515;
        else
            _1516 <= _1513;
    end
    always @(posedge _84) begin
        if (_82)
            _1519 <= _1518;
        else
            _1519 <= _1516;
    end
    always @(posedge _84) begin
        if (_82)
            _1522 <= _1521;
        else
            _1522 <= _1519;
    end
    always @(posedge _84) begin
        if (_82)
            _1525 <= _1524;
        else
            _1525 <= _1522;
    end
    always @(posedge _84) begin
        if (_82)
            _1528 <= _1527;
        else
            _1528 <= _1525;
    end
    always @(posedge _84) begin
        if (_82)
            _1531 <= _1530;
        else
            _1531 <= _1528;
    end
    assign _1532 = ~ _1531;
    always @(posedge _84) begin
        if (_82)
            _1480 <= _1479;
        else
            _1480 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1483 <= _1482;
        else
            _1483 <= _1480;
    end
    always @(posedge _84) begin
        if (_82)
            _1486 <= _1485;
        else
            _1486 <= _1483;
    end
    always @(posedge _84) begin
        if (_82)
            _1489 <= _1488;
        else
            _1489 <= _1486;
    end
    always @(posedge _84) begin
        if (_82)
            _1492 <= _1491;
        else
            _1492 <= _1489;
    end
    always @(posedge _84) begin
        if (_82)
            _1495 <= _1494;
        else
            _1495 <= _1492;
    end
    always @(posedge _84) begin
        if (_82)
            _1498 <= _1497;
        else
            _1498 <= _1495;
    end
    always @(posedge _84) begin
        if (_82)
            _1501 <= _1500;
        else
            _1501 <= _1498;
    end
    always @(posedge _84) begin
        if (_82)
            _1504 <= _1503;
        else
            _1504 <= _1501;
    end
    assign _1533 = _1504 & _1532;
    assign _1534 = _129 & _1533;
    assign write_enable_82 = _1534 & PHASE_19;
    assign _1539 = write_enable_82 | read_enable_68;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_40
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1539), .regcea(vdd), .wea(write_enable_82), .addra(address_82), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_73), .regceb(vdd), .web(write_enable_73), .addrb(address_73), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1546[131:131]), .sbiterrb(_1546[130:130]), .doutb(_1546[129:66]), .dbiterra(_1546[65:65]), .sbiterra(_1546[64:64]), .douta(_1546[63:0]) );
    assign _1547 = _1546[63:0];
    assign _1477 = ~ PHASE_19;
    assign _55 = _1477;
    always @(posedge _84) begin
        if (_82)
            PHASE_19 <= _1475;
        else
            if (_72)
                PHASE_19 <= _55;
    end
    assign _1559 = PHASE_19 ? _1558 : _1547;
    assign address_83 = _1744 ? _199 : _1739;
    assign write_enable_83 = _1737 & _1744;
    assign address_84 = _1744 ? _164 : _68;
    assign _1746 = ~ _1744;
    assign read_enable_69 = _1732 & _1746;
    assign _1744 = ~ PHASE_22;
    assign write_enable_84 = _1730 & _1744;
    assign _1748 = write_enable_84 | read_enable_69;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_41
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1748), .regcea(vdd), .wea(write_enable_84), .addra(address_84), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_83), .regceb(vdd), .web(write_enable_83), .addrb(address_83), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1753[131:131]), .sbiterrb(_1753[130:130]), .doutb(_1753[129:66]), .dbiterra(_1753[65:65]), .sbiterra(_1753[64:64]), .douta(_1753[63:0]) );
    assign _1754 = _1753[63:0];
    assign address_85 = PHASE_22 ? _199 : _1739;
    assign _1737 = _129 & _1700;
    assign write_enable_85 = _1737 & PHASE_22;
    assign _292 = _91[521:518];
    assign _291 = _91[517:517];
    assign _289 = _91[513:513];
    assign _288 = _91[512:449];
    assign _287 = _91[448:385];
    assign _286 = _91[384:321];
    assign _285 = _91[320:257];
    assign _284 = _91[256:193];
    assign _283 = _91[192:129];
    assign _282 = _91[128:65];
    assign _1662 = _1654[129:66];
    assign _1661 = _1641[129:66];
    assign _1663 = PHASE_20 ? _1662 : _1661;
    assign _1659 = _1599[129:66];
    assign _1658 = _1585[129:66];
    assign q1_6 = PHASE_21 ? _1659 : _1658;
    assign _1664 = _1566 ? _1663 : q1_6;
    assign address_86 = _1643 ? _1637 : _1636;
    assign _1649 = ~ _1643;
    assign read_enable_70 = _102 & _1649;
    assign address_87 = _1643 ? _60 : _1619;
    assign _1645 = ~ _1643;
    assign read_enable_71 = _102 & _1645;
    assign _1643 = ~ PHASE_20;
    assign write_enable_87 = _1602 & _1643;
    assign _1647 = write_enable_87 | read_enable_71;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_42
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1647), .regcea(vdd), .wea(write_enable_87), .addra(address_87), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_70), .regceb(vdd), .web(write_enable_86), .addrb(address_86), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1654[131:131]), .sbiterrb(_1654[130:130]), .doutb(_1654[129:66]), .dbiterra(_1654[65:65]), .sbiterra(_1654[64:64]), .douta(_1654[63:0]) );
    assign _1655 = _1654[63:0];
    assign _1635 = _172[11:11];
    assign _1634 = _172[10:10];
    assign _1633 = _172[9:9];
    assign _1632 = _172[8:8];
    assign _1631 = _172[7:7];
    assign _1630 = _172[6:6];
    assign _1629 = _172[5:5];
    assign _1628 = _172[4:4];
    assign _1627 = _172[3:3];
    assign _1626 = _172[2:2];
    assign _1625 = _172[1:1];
    assign _1624 = _172[0:0];
    assign _1636 = { _1624, _1625, _1626, _1627, _1628, _1629, _1630, _1631, _1632, _1633, _1634, _1635 };
    assign address_88 = PHASE_20 ? _1637 : _1636;
    assign _1621 = ~ PHASE_20;
    assign read_enable_72 = _102 & _1621;
    assign data_85 = wr_d0;
    assign _60 = wr_addr;
    assign _1618 = _137[11:11];
    assign _1617 = _137[10:10];
    assign _1616 = _137[9:9];
    assign _1615 = _137[8:8];
    assign _1614 = _137[7:7];
    assign _1613 = _137[6:6];
    assign _1612 = _137[5:5];
    assign _1611 = _137[4:4];
    assign _1610 = _137[3:3];
    assign _1609 = _137[2:2];
    assign _1608 = _137[1:1];
    assign _1607 = _137[0:0];
    assign _1619 = { _1607, _1608, _1609, _1610, _1611, _1612, _1613, _1614, _1615, _1616, _1617, _1618 };
    assign address_89 = PHASE_20 ? _60 : _1619;
    assign _1604 = ~ PHASE_20;
    assign read_enable_73 = _102 & _1604;
    assign _62 = wr_en;
    assign _1602 = _62[0:0];
    assign write_enable_89 = _1602 & PHASE_20;
    assign _1606 = write_enable_89 | read_enable_73;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_43
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1606), .regcea(vdd), .wea(write_enable_89), .addra(address_89), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_72), .regceb(vdd), .web(write_enable_88), .addrb(address_88), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1641[131:131]), .sbiterrb(_1641[130:130]), .doutb(_1641[129:66]), .dbiterra(_1641[65:65]), .sbiterra(_1641[64:64]), .douta(_1641[63:0]) );
    assign _1642 = _1641[63:0];
    assign _1563 = ~ PHASE_20;
    assign _63 = _1563;
    always @(posedge _84) begin
        if (_82)
            PHASE_20 <= _1561;
        else
            if (_72)
                PHASE_20 <= _63;
    end
    assign _1656 = PHASE_20 ? _1655 : _1642;
    assign address_90 = _1587 ? _199 : _172;
    assign _1594 = ~ _1587;
    assign read_enable_74 = _102 & _1594;
    assign write_enable_90 = _1578 & _1587;
    assign _1596 = write_enable_90 | read_enable_74;
    assign address_91 = _1587 ? _164 : _137;
    assign _1589 = ~ _1587;
    assign read_enable_75 = _102 & _1589;
    assign _1587 = ~ PHASE_21;
    assign write_enable_91 = _1571 & _1587;
    assign _1591 = write_enable_91 | read_enable_75;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_44
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1591), .regcea(vdd), .wea(write_enable_91), .addra(address_91), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1596), .regceb(vdd), .web(write_enable_90), .addrb(address_90), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1599[131:131]), .sbiterrb(_1599[130:130]), .doutb(_1599[129:66]), .dbiterra(_1599[65:65]), .sbiterra(_1599[64:64]), .douta(_1599[63:0]) );
    assign _1600 = _1599[63:0];
    assign _1667 = _1666[127:64];
    assign data_87 = _1667;
    always @(posedge _84) begin
        if (_82)
            _175 <= _174;
        else
            _175 <= _172;
    end
    always @(posedge _84) begin
        if (_82)
            _178 <= _177;
        else
            _178 <= _175;
    end
    always @(posedge _84) begin
        if (_82)
            _181 <= _180;
        else
            _181 <= _178;
    end
    always @(posedge _84) begin
        if (_82)
            _184 <= _183;
        else
            _184 <= _181;
    end
    always @(posedge _84) begin
        if (_82)
            _187 <= _186;
        else
            _187 <= _184;
    end
    always @(posedge _84) begin
        if (_82)
            _190 <= _189;
        else
            _190 <= _187;
    end
    always @(posedge _84) begin
        if (_82)
            _193 <= _192;
        else
            _193 <= _190;
    end
    always @(posedge _84) begin
        if (_82)
            _196 <= _195;
        else
            _196 <= _193;
    end
    always @(posedge _84) begin
        if (_82)
            _199 <= _198;
        else
            _199 <= _196;
    end
    assign _172 = _91[64:53];
    assign address_92 = PHASE_21 ? _199 : _172;
    assign _1580 = ~ PHASE_21;
    assign read_enable_76 = _102 & _1580;
    assign _1577 = ~ _130;
    assign _1578 = _129 & _1577;
    assign write_enable_92 = _1578 & PHASE_21;
    assign _1582 = write_enable_92 | read_enable_76;
    assign address_93 = PHASE_21 ? _164 : _137;
    assign _1573 = ~ PHASE_21;
    assign read_enable_77 = _102 & _1573;
    assign _1570 = ~ _130;
    assign _1571 = _129 & _1570;
    assign write_enable_93 = _1571 & PHASE_21;
    assign _1575 = write_enable_93 | read_enable_77;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_45
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1575), .regcea(vdd), .wea(write_enable_93), .addra(address_93), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1582), .regceb(vdd), .web(write_enable_92), .addrb(address_92), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1585[131:131]), .sbiterrb(_1585[130:130]), .doutb(_1585[129:66]), .dbiterra(_1585[65:65]), .sbiterra(_1585[64:64]), .douta(_1585[63:0]) );
    assign _1586 = _1585[63:0];
    assign _99 = _91[523:523];
    assign _1668 = ~ PHASE_21;
    assign _65 = _1668;
    always @(posedge _84) begin
        if (_82)
            PHASE_21 <= _1568;
        else
            if (_99)
                PHASE_21 <= _65;
    end
    assign q0_6 = PHASE_21 ? _1600 : _1586;
    assign _92 = _91[514:514];
    always @(posedge _84) begin
        if (_82)
            _1566 <= _1565;
        else
            _1566 <= _92;
    end
    assign _1657 = _1566 ? _1656 : q0_6;
    dp_39
        dp
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1657), .d2(_1664), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1666[191:128]), .q2(_1666[127:64]), .q1(_1666[63:0]) );
    assign _1669 = _1666[63:0];
    assign data_91 = _1669;
    assign _137 = _91[52:41];
    always @(posedge _84) begin
        if (_82)
            _140 <= _139;
        else
            _140 <= _137;
    end
    always @(posedge _84) begin
        if (_82)
            _143 <= _142;
        else
            _143 <= _140;
    end
    always @(posedge _84) begin
        if (_82)
            _146 <= _145;
        else
            _146 <= _143;
    end
    always @(posedge _84) begin
        if (_82)
            _149 <= _148;
        else
            _149 <= _146;
    end
    always @(posedge _84) begin
        if (_82)
            _152 <= _151;
        else
            _152 <= _149;
    end
    always @(posedge _84) begin
        if (_82)
            _155 <= _154;
        else
            _155 <= _152;
    end
    always @(posedge _84) begin
        if (_82)
            _158 <= _157;
        else
            _158 <= _155;
    end
    always @(posedge _84) begin
        if (_82)
            _161 <= _160;
        else
            _161 <= _158;
    end
    always @(posedge _84) begin
        if (_82)
            _164 <= _163;
        else
            _164 <= _161;
    end
    assign _68 = rd_addr;
    assign address_94 = PHASE_22 ? _164 : _68;
    assign _1733 = ~ PHASE_22;
    assign _70 = rd_en;
    assign _1732 = _70[0:0];
    assign read_enable_78 = _1732 & _1733;
    assign _290 = _91[516:516];
    always @(posedge _84) begin
        if (_82)
            _1703 <= _1702;
        else
            _1703 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1706 <= _1705;
        else
            _1706 <= _1703;
    end
    always @(posedge _84) begin
        if (_82)
            _1709 <= _1708;
        else
            _1709 <= _1706;
    end
    always @(posedge _84) begin
        if (_82)
            _1712 <= _1711;
        else
            _1712 <= _1709;
    end
    always @(posedge _84) begin
        if (_82)
            _1715 <= _1714;
        else
            _1715 <= _1712;
    end
    always @(posedge _84) begin
        if (_82)
            _1718 <= _1717;
        else
            _1718 <= _1715;
    end
    always @(posedge _84) begin
        if (_82)
            _1721 <= _1720;
        else
            _1721 <= _1718;
    end
    always @(posedge _84) begin
        if (_82)
            _1724 <= _1723;
        else
            _1724 <= _1721;
    end
    always @(posedge _84) begin
        if (_82)
            _1727 <= _1726;
        else
            _1727 <= _1724;
    end
    assign _1728 = ~ _1727;
    assign _130 = _91[515:515];
    always @(posedge _84) begin
        if (_82)
            _1676 <= _1675;
        else
            _1676 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1679 <= _1678;
        else
            _1679 <= _1676;
    end
    always @(posedge _84) begin
        if (_82)
            _1682 <= _1681;
        else
            _1682 <= _1679;
    end
    always @(posedge _84) begin
        if (_82)
            _1685 <= _1684;
        else
            _1685 <= _1682;
    end
    always @(posedge _84) begin
        if (_82)
            _1688 <= _1687;
        else
            _1688 <= _1685;
    end
    always @(posedge _84) begin
        if (_82)
            _1691 <= _1690;
        else
            _1691 <= _1688;
    end
    always @(posedge _84) begin
        if (_82)
            _1694 <= _1693;
        else
            _1694 <= _1691;
    end
    always @(posedge _84) begin
        if (_82)
            _1697 <= _1696;
        else
            _1697 <= _1694;
    end
    always @(posedge _84) begin
        if (_82)
            _1700 <= _1699;
        else
            _1700 <= _1697;
    end
    assign _1729 = _1700 & _1728;
    assign _102 = _91[522:522];
    always @(posedge _84) begin
        if (_82)
            _105 <= _104;
        else
            _105 <= _102;
    end
    always @(posedge _84) begin
        if (_82)
            _108 <= _107;
        else
            _108 <= _105;
    end
    always @(posedge _84) begin
        if (_82)
            _111 <= _110;
        else
            _111 <= _108;
    end
    always @(posedge _84) begin
        if (_82)
            _114 <= _113;
        else
            _114 <= _111;
    end
    always @(posedge _84) begin
        if (_82)
            _117 <= _116;
        else
            _117 <= _114;
    end
    always @(posedge _84) begin
        if (_82)
            _120 <= _119;
        else
            _120 <= _117;
    end
    always @(posedge _84) begin
        if (_82)
            _123 <= _122;
        else
            _123 <= _120;
    end
    always @(posedge _84) begin
        if (_82)
            _126 <= _125;
        else
            _126 <= _123;
    end
    always @(posedge _84) begin
        if (_82)
            _129 <= _128;
        else
            _129 <= _126;
    end
    assign _1730 = _129 & _1729;
    assign write_enable_94 = _1730 & PHASE_22;
    assign _1735 = write_enable_94 | read_enable_78;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_46
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1735), .regcea(vdd), .wea(write_enable_94), .addra(address_94), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_85), .regceb(vdd), .web(write_enable_85), .addrb(address_85), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1742[131:131]), .sbiterrb(_1742[130:130]), .doutb(_1742[129:66]), .dbiterra(_1742[65:65]), .sbiterra(_1742[64:64]), .douta(_1742[63:0]) );
    assign _1743 = _1742[63:0];
    assign _72 = flip;
    assign _1673 = ~ PHASE_22;
    assign _73 = _1673;
    always @(posedge _84) begin
        if (_82)
            PHASE_22 <= _1671;
        else
            if (_72)
                PHASE_22 <= _73;
    end
    assign _1755 = PHASE_22 ? _1754 : _1743;
    assign _76 = first_4step_pass;
    assign _78 = first_iter;
    assign _80 = start;
    assign _82 = clear;
    assign _84 = clock;
    ctrl
        ctrl
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .first_4step_pass(_76), .flip(_91[523:523]), .read_write_enable(_91[522:522]), .index(_91[521:518]), .valid(_91[517:517]), .twiddle_stage(_91[516:516]), .last_stage(_91[515:515]), .first_stage(_91[514:514]), .start_twiddles(_91[513:513]), .omegas6(_91[512:449]), .omegas5(_91[448:385]), .omegas4(_91[384:321]), .omegas3(_91[320:257]), .omegas2(_91[256:193]), .omegas1(_91[192:129]), .omegas0(_91[128:65]), .addr2(_91[64:53]), .addr1(_91[52:41]), .m(_91[40:29]), .k(_91[28:17]), .j(_91[16:5]), .i(_91[4:1]), .done_(_91[0:0]) );
    assign _1756 = _91[0:0];

    /* aliases */
    assign data_0 = data;
    assign data_2 = data_1;
    assign data_4 = data_3;
    assign data_5 = data_3;
    assign data_6 = data_3;
    assign data_8 = data_7;
    assign data_9 = data_7;
    assign data_10 = data_7;
    assign data_12 = data_11;
    assign data_14 = data_13;
    assign data_16 = data_15;
    assign data_17 = data_15;
    assign data_18 = data_15;
    assign data_20 = data_19;
    assign data_21 = data_19;
    assign data_22 = data_19;
    assign data_24 = data_23;
    assign data_26 = data_25;
    assign data_28 = data_27;
    assign data_29 = data_27;
    assign data_30 = data_27;
    assign data_32 = data_31;
    assign data_33 = data_31;
    assign data_34 = data_31;
    assign data_36 = data_35;
    assign data_38 = data_37;
    assign data_40 = data_39;
    assign data_41 = data_39;
    assign data_42 = data_39;
    assign data_44 = data_43;
    assign data_45 = data_43;
    assign data_46 = data_43;
    assign data_48 = data_47;
    assign data_50 = data_49;
    assign data_52 = data_51;
    assign data_53 = data_51;
    assign data_54 = data_51;
    assign data_56 = data_55;
    assign data_57 = data_55;
    assign data_58 = data_55;
    assign data_60 = data_59;
    assign data_62 = data_61;
    assign data_64 = data_63;
    assign data_65 = data_63;
    assign data_66 = data_63;
    assign data_68 = data_67;
    assign data_69 = data_67;
    assign data_70 = data_67;
    assign data_72 = data_71;
    assign data_74 = data_73;
    assign data_76 = data_75;
    assign data_77 = data_75;
    assign data_78 = data_75;
    assign data_80 = data_79;
    assign data_81 = data_79;
    assign data_82 = data_79;
    assign data_84 = data_83;
    assign data_86 = data_85;
    assign data_88 = data_87;
    assign data_89 = data_87;
    assign data_90 = data_87;
    assign data_92 = data_91;
    assign data_93 = data_91;
    assign data_94 = data_91;

    /* output assignments */
    assign done_ = _1756;
    assign rd_q0 = _1755;
    assign rd_q1 = _1559;
    assign rd_q2 = _1363;
    assign rd_q3 = _1167;
    assign rd_q4 = _971;
    assign rd_q5 = _775;
    assign rd_q6 = _579;
    assign rd_q7 = _383;

endmodule
module dp_47 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1011110000101000110110001111100101001011011110101100100100000000;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0001011100110100000001011010010010001110111001001000001101001101;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0000010100000011100011000110011101011000001110100111010001011001;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0011110101010110000000001101011100010100100101111100001010111100;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0110100110010111111010001101100011001001101111010100100000100101;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0000101011001010001100100100101101011011001100100000011011011100;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_48 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1010100110000001001000000000101010100000110110001011101001110101;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0000101110000011010000000101110111010110101101011011110001111001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1101011010101010101100111101101011101110011110100000110011000011;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1001001111001111100100101110011001000010100110100100110010010011;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0101000011001111001101110000000110110101011011100101101000110110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1000000110101110110111001110001000000110110000010101010010110101;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0010100101000101111001010011010000000110010111011010001100101101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_49 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0111111100000111000101010111111111111011100111110111010001111100;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0110011000111100001011010000011010111111001001111000111011100101;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1010101101110001111011100110111011001110000111110011100011101010;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0001011001000100000110101011001011011010101100111100000011000001;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1000101101111010111110100101101000010010011111110000010100011000;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0001011111010001110111110010100111110100110100010110100100111010;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0001100100000101011100000100110001000100110010001101110010111010;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_50 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0101101110010110010100001111010010111110001000010100011011111011;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1000001001111101111011000100111100101011100011100001010111001110;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0001100110101110101010110011101100000101001000111001100000000011;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0000101111001000100000001011001110110011001101111111011010000101;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0110110001110101010111000111101110001101010111001100011001010000;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0111111010110111000101110011011011100010101100111010000100000110;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0110000010001000010110101101110010000100111001101000101001111110;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_51 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1000100110110001111010000001100001011111100010101001100011001100;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0100110010001001010001111001010000110110101011101010001000000001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1000111001000111011111010100101000111011010001000110101100010010;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0011111111100110010011010010011110110101100101011111011101111100;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0110101010010110110001001110100010101101100101010001110111001100;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0110010010111101011010101001111010001000110111100110011111100000;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1000011011100101001000010011100100111101111001011101100010110100;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_52 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0111010100011100101000100011001111101000111010111111001001111101;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1011010110111101100001101100000111110001011001011001110000010000;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0101111110110010100111011111111111111110011010100111101111101100;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0010110110111110111001110010010110100101000011101110000110100010;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0111101100101101010001110010010110001011011001100000111110111000;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1010011011000111110110011110001000111001000110110100110011010000;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1001001000110110001100101001101010110111011101111111000111011010;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_53 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0011011011110011000011111101110100101011011111110100100011001001;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1100111011001100001100110110110100110010010011010100111111001011;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1111000101010111111011100011110110011011001000100001010100111100;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b1010001101101010010111100101011111010001100010010100010001010001;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1111101101011111000100111011001000110101001100000101010001101001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0001001000111000010111110001101011011001000001111111010110000000;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0000000010100111001011000000010010100111011101011111110001111000;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_54 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0100011011000000110111000111111100101001111000011000110101111010;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0000101111110001010101001100101001111110111001110111010001010000;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0101101000000110010100101010000011101000100001011010011110010001;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0010000101110010001101000110101010000001001100100101001010100011;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0100001010110000001101000000101010000000011110111001101000111101;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1001010100101001000110000101000110101101100000000110001101010110;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0000110011111011010001010110001011100101111101011000011111100101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module parallel_cores_5 (
    wr_d7,
    wr_d6,
    wr_d5,
    wr_d4,
    wr_d3,
    wr_d2,
    wr_d1,
    wr_d0,
    wr_addr,
    wr_en,
    rd_addr,
    rd_en,
    flip,
    first_4step_pass,
    first_iter,
    start,
    clear,
    clock,
    done_,
    rd_q0,
    rd_q1,
    rd_q2,
    rd_q3,
    rd_q4,
    rd_q5,
    rd_q6,
    rd_q7
);

    input [63:0] wr_d7;
    input [63:0] wr_d6;
    input [63:0] wr_d5;
    input [63:0] wr_d4;
    input [63:0] wr_d3;
    input [63:0] wr_d2;
    input [63:0] wr_d1;
    input [63:0] wr_d0;
    input [11:0] wr_addr;
    input [7:0] wr_en;
    input [11:0] rd_addr;
    input [7:0] rd_en;
    input flip;
    input first_4step_pass;
    input first_iter;
    input start;
    input clear;
    input clock;
    output done_;
    output [63:0] rd_q0;
    output [63:0] rd_q1;
    output [63:0] rd_q2;
    output [63:0] rd_q3;
    output [63:0] rd_q4;
    output [63:0] rd_q5;
    output [63:0] rd_q6;
    output [63:0] rd_q7;

    /* signal declarations */
    wire [11:0] address;
    wire write_enable;
    wire [11:0] address_0;
    wire _374;
    wire read_enable;
    wire _372;
    wire write_enable_0;
    wire _376;
    wire [131:0] _381;
    wire [63:0] _382;
    wire [11:0] _367 = 12'b000000000000;
    wire [11:0] address_1;
    wire _365;
    wire write_enable_1;
    wire [63:0] _279;
    wire [63:0] _278;
    wire [63:0] _280;
    wire [63:0] _276;
    wire [63:0] _275;
    wire [63:0] q1;
    wire [63:0] _281;
    wire [11:0] address_2;
    wire write_enable_2 = 1'b0;
    wire _266;
    wire read_enable_0;
    wire [11:0] address_3;
    wire _262;
    wire read_enable_1;
    wire _260;
    wire write_enable_3;
    wire _264;
    wire [131:0] _271;
    wire [63:0] _272;
    wire [63:0] data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_0;
    wire [11:0] _254 = 12'b000000000000;
    wire _252;
    wire _251;
    wire _250;
    wire _249;
    wire _248;
    wire _247;
    wire _246;
    wire _245;
    wire _244;
    wire _243;
    wire _242;
    wire _241;
    wire [11:0] _253;
    wire [11:0] address_4;
    wire write_enable_4 = 1'b0;
    wire _238;
    wire read_enable_2;
    wire [63:0] data_1;
    wire [63:0] data_2;
    wire _235;
    wire _234;
    wire _233;
    wire _232;
    wire _231;
    wire _230;
    wire _229;
    wire _228;
    wire _227;
    wire _226;
    wire _225;
    wire _224;
    wire [11:0] _236;
    wire [11:0] address_5;
    wire _221;
    wire read_enable_3;
    wire _219;
    wire write_enable_5;
    wire _223;
    wire [131:0] _258;
    wire [63:0] _259;
    wire _87 = 1'b0;
    wire _86 = 1'b0;
    wire _89;
    wire _3;
    reg PHASE;
    wire [63:0] _273;
    wire [11:0] address_6;
    wire _211;
    wire read_enable_4;
    wire write_enable_6;
    wire _213;
    wire [11:0] address_7;
    wire _206;
    wire read_enable_5;
    wire _204;
    wire write_enable_7;
    wire _208;
    wire [131:0] _216;
    wire [63:0] _217;
    wire [63:0] _295;
    wire [63:0] data_3;
    wire [63:0] data_4;
    wire [63:0] data_5;
    wire [63:0] data_6;
    wire [11:0] address_8;
    wire _169;
    wire read_enable_6;
    wire _166;
    wire _167;
    wire write_enable_8;
    wire _171;
    wire [11:0] address_9;
    wire _134;
    wire read_enable_7;
    wire _131;
    wire _132;
    wire write_enable_9;
    wire _136;
    wire [131:0] _202;
    wire [63:0] _203;
    wire _98 = 1'b0;
    wire _97 = 1'b0;
    wire _296;
    wire _5;
    reg PHASE_0;
    wire [63:0] q0;
    wire _94 = 1'b0;
    wire _93 = 1'b0;
    reg _96;
    wire [63:0] _274;
    wire [191:0] _294;
    wire [63:0] _297;
    wire [63:0] data_7;
    wire [63:0] data_8;
    wire [63:0] data_9;
    wire [63:0] data_10;
    wire [11:0] address_10;
    wire _361;
    wire _360;
    wire read_enable_8;
    wire _354 = 1'b0;
    wire _353 = 1'b0;
    wire _351 = 1'b0;
    wire _350 = 1'b0;
    wire _348 = 1'b0;
    wire _347 = 1'b0;
    wire _345 = 1'b0;
    wire _344 = 1'b0;
    wire _342 = 1'b0;
    wire _341 = 1'b0;
    wire _339 = 1'b0;
    wire _338 = 1'b0;
    wire _336 = 1'b0;
    wire _335 = 1'b0;
    wire _333 = 1'b0;
    wire _332 = 1'b0;
    wire _330 = 1'b0;
    wire _329 = 1'b0;
    reg _331;
    reg _334;
    reg _337;
    reg _340;
    reg _343;
    reg _346;
    reg _349;
    reg _352;
    reg _355;
    wire _356;
    wire _327 = 1'b0;
    wire _326 = 1'b0;
    wire _324 = 1'b0;
    wire _323 = 1'b0;
    wire _321 = 1'b0;
    wire _320 = 1'b0;
    wire _318 = 1'b0;
    wire _317 = 1'b0;
    wire _315 = 1'b0;
    wire _314 = 1'b0;
    wire _312 = 1'b0;
    wire _311 = 1'b0;
    wire _309 = 1'b0;
    wire _308 = 1'b0;
    wire _306 = 1'b0;
    wire _305 = 1'b0;
    wire _303 = 1'b0;
    wire _302 = 1'b0;
    reg _304;
    reg _307;
    reg _310;
    reg _313;
    reg _316;
    reg _319;
    reg _322;
    reg _325;
    reg _328;
    wire _357;
    wire _358;
    wire write_enable_10;
    wire _363;
    wire [131:0] _370;
    wire [63:0] _371;
    wire _299 = 1'b0;
    wire _298 = 1'b0;
    wire _301;
    wire _7;
    reg PHASE_1;
    wire [63:0] _383;
    wire [11:0] address_11;
    wire write_enable_11;
    wire [11:0] address_12;
    wire _570;
    wire read_enable_9;
    wire _568;
    wire write_enable_12;
    wire _572;
    wire [131:0] _577;
    wire [63:0] _578;
    wire [11:0] _563 = 12'b000000000000;
    wire [11:0] address_13;
    wire _561;
    wire write_enable_13;
    wire [63:0] _486;
    wire [63:0] _485;
    wire [63:0] _487;
    wire [63:0] _483;
    wire [63:0] _482;
    wire [63:0] q1_0;
    wire [63:0] _488;
    wire [11:0] address_14;
    wire write_enable_14 = 1'b0;
    wire _473;
    wire read_enable_10;
    wire [11:0] address_15;
    wire _469;
    wire read_enable_11;
    wire _467;
    wire write_enable_15;
    wire _471;
    wire [131:0] _478;
    wire [63:0] _479;
    wire [63:0] data_11 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_12;
    wire [11:0] _461 = 12'b000000000000;
    wire _459;
    wire _458;
    wire _457;
    wire _456;
    wire _455;
    wire _454;
    wire _453;
    wire _452;
    wire _451;
    wire _450;
    wire _449;
    wire _448;
    wire [11:0] _460;
    wire [11:0] address_16;
    wire write_enable_16 = 1'b0;
    wire _445;
    wire read_enable_12;
    wire [63:0] data_13;
    wire [63:0] data_14;
    wire _442;
    wire _441;
    wire _440;
    wire _439;
    wire _438;
    wire _437;
    wire _436;
    wire _435;
    wire _434;
    wire _433;
    wire _432;
    wire _431;
    wire [11:0] _443;
    wire [11:0] address_17;
    wire _428;
    wire read_enable_13;
    wire _426;
    wire write_enable_17;
    wire _430;
    wire [131:0] _465;
    wire [63:0] _466;
    wire _385 = 1'b0;
    wire _384 = 1'b0;
    wire _387;
    wire _11;
    reg PHASE_2;
    wire [63:0] _480;
    wire [11:0] address_18;
    wire _418;
    wire read_enable_14;
    wire write_enable_18;
    wire _420;
    wire [11:0] address_19;
    wire _413;
    wire read_enable_15;
    wire _411;
    wire write_enable_19;
    wire _415;
    wire [131:0] _423;
    wire [63:0] _424;
    wire [63:0] _491;
    wire [63:0] data_15;
    wire [63:0] data_16;
    wire [63:0] data_17;
    wire [63:0] data_18;
    wire [11:0] address_20;
    wire _404;
    wire read_enable_16;
    wire _401;
    wire _402;
    wire write_enable_20;
    wire _406;
    wire [11:0] address_21;
    wire _397;
    wire read_enable_17;
    wire _394;
    wire _395;
    wire write_enable_21;
    wire _399;
    wire [131:0] _409;
    wire [63:0] _410;
    wire _392 = 1'b0;
    wire _391 = 1'b0;
    wire _492;
    wire _13;
    reg PHASE_3;
    wire [63:0] q0_0;
    wire _389 = 1'b0;
    wire _388 = 1'b0;
    reg _390;
    wire [63:0] _481;
    wire [191:0] _490;
    wire [63:0] _493;
    wire [63:0] data_19;
    wire [63:0] data_20;
    wire [63:0] data_21;
    wire [63:0] data_22;
    wire [11:0] address_22;
    wire _557;
    wire _556;
    wire read_enable_18;
    wire _550 = 1'b0;
    wire _549 = 1'b0;
    wire _547 = 1'b0;
    wire _546 = 1'b0;
    wire _544 = 1'b0;
    wire _543 = 1'b0;
    wire _541 = 1'b0;
    wire _540 = 1'b0;
    wire _538 = 1'b0;
    wire _537 = 1'b0;
    wire _535 = 1'b0;
    wire _534 = 1'b0;
    wire _532 = 1'b0;
    wire _531 = 1'b0;
    wire _529 = 1'b0;
    wire _528 = 1'b0;
    wire _526 = 1'b0;
    wire _525 = 1'b0;
    reg _527;
    reg _530;
    reg _533;
    reg _536;
    reg _539;
    reg _542;
    reg _545;
    reg _548;
    reg _551;
    wire _552;
    wire _523 = 1'b0;
    wire _522 = 1'b0;
    wire _520 = 1'b0;
    wire _519 = 1'b0;
    wire _517 = 1'b0;
    wire _516 = 1'b0;
    wire _514 = 1'b0;
    wire _513 = 1'b0;
    wire _511 = 1'b0;
    wire _510 = 1'b0;
    wire _508 = 1'b0;
    wire _507 = 1'b0;
    wire _505 = 1'b0;
    wire _504 = 1'b0;
    wire _502 = 1'b0;
    wire _501 = 1'b0;
    wire _499 = 1'b0;
    wire _498 = 1'b0;
    reg _500;
    reg _503;
    reg _506;
    reg _509;
    reg _512;
    reg _515;
    reg _518;
    reg _521;
    reg _524;
    wire _553;
    wire _554;
    wire write_enable_22;
    wire _559;
    wire [131:0] _566;
    wire [63:0] _567;
    wire _495 = 1'b0;
    wire _494 = 1'b0;
    wire _497;
    wire _15;
    reg PHASE_4;
    wire [63:0] _579;
    wire [11:0] address_23;
    wire write_enable_23;
    wire [11:0] address_24;
    wire _766;
    wire read_enable_19;
    wire _764;
    wire write_enable_24;
    wire _768;
    wire [131:0] _773;
    wire [63:0] _774;
    wire [11:0] _759 = 12'b000000000000;
    wire [11:0] address_25;
    wire _757;
    wire write_enable_25;
    wire [63:0] _682;
    wire [63:0] _681;
    wire [63:0] _683;
    wire [63:0] _679;
    wire [63:0] _678;
    wire [63:0] q1_1;
    wire [63:0] _684;
    wire [11:0] address_26;
    wire write_enable_26 = 1'b0;
    wire _669;
    wire read_enable_20;
    wire [11:0] address_27;
    wire _665;
    wire read_enable_21;
    wire _663;
    wire write_enable_27;
    wire _667;
    wire [131:0] _674;
    wire [63:0] _675;
    wire [63:0] data_23 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_24;
    wire [11:0] _657 = 12'b000000000000;
    wire _655;
    wire _654;
    wire _653;
    wire _652;
    wire _651;
    wire _650;
    wire _649;
    wire _648;
    wire _647;
    wire _646;
    wire _645;
    wire _644;
    wire [11:0] _656;
    wire [11:0] address_28;
    wire write_enable_28 = 1'b0;
    wire _641;
    wire read_enable_22;
    wire [63:0] data_25;
    wire [63:0] data_26;
    wire _638;
    wire _637;
    wire _636;
    wire _635;
    wire _634;
    wire _633;
    wire _632;
    wire _631;
    wire _630;
    wire _629;
    wire _628;
    wire _627;
    wire [11:0] _639;
    wire [11:0] address_29;
    wire _624;
    wire read_enable_23;
    wire _622;
    wire write_enable_29;
    wire _626;
    wire [131:0] _661;
    wire [63:0] _662;
    wire _581 = 1'b0;
    wire _580 = 1'b0;
    wire _583;
    wire _19;
    reg PHASE_5;
    wire [63:0] _676;
    wire [11:0] address_30;
    wire _614;
    wire read_enable_24;
    wire write_enable_30;
    wire _616;
    wire [11:0] address_31;
    wire _609;
    wire read_enable_25;
    wire _607;
    wire write_enable_31;
    wire _611;
    wire [131:0] _619;
    wire [63:0] _620;
    wire [63:0] _687;
    wire [63:0] data_27;
    wire [63:0] data_28;
    wire [63:0] data_29;
    wire [63:0] data_30;
    wire [11:0] address_32;
    wire _600;
    wire read_enable_26;
    wire _597;
    wire _598;
    wire write_enable_32;
    wire _602;
    wire [11:0] address_33;
    wire _593;
    wire read_enable_27;
    wire _590;
    wire _591;
    wire write_enable_33;
    wire _595;
    wire [131:0] _605;
    wire [63:0] _606;
    wire _588 = 1'b0;
    wire _587 = 1'b0;
    wire _688;
    wire _21;
    reg PHASE_6;
    wire [63:0] q0_1;
    wire _585 = 1'b0;
    wire _584 = 1'b0;
    reg _586;
    wire [63:0] _677;
    wire [191:0] _686;
    wire [63:0] _689;
    wire [63:0] data_31;
    wire [63:0] data_32;
    wire [63:0] data_33;
    wire [63:0] data_34;
    wire [11:0] address_34;
    wire _753;
    wire _752;
    wire read_enable_28;
    wire _746 = 1'b0;
    wire _745 = 1'b0;
    wire _743 = 1'b0;
    wire _742 = 1'b0;
    wire _740 = 1'b0;
    wire _739 = 1'b0;
    wire _737 = 1'b0;
    wire _736 = 1'b0;
    wire _734 = 1'b0;
    wire _733 = 1'b0;
    wire _731 = 1'b0;
    wire _730 = 1'b0;
    wire _728 = 1'b0;
    wire _727 = 1'b0;
    wire _725 = 1'b0;
    wire _724 = 1'b0;
    wire _722 = 1'b0;
    wire _721 = 1'b0;
    reg _723;
    reg _726;
    reg _729;
    reg _732;
    reg _735;
    reg _738;
    reg _741;
    reg _744;
    reg _747;
    wire _748;
    wire _719 = 1'b0;
    wire _718 = 1'b0;
    wire _716 = 1'b0;
    wire _715 = 1'b0;
    wire _713 = 1'b0;
    wire _712 = 1'b0;
    wire _710 = 1'b0;
    wire _709 = 1'b0;
    wire _707 = 1'b0;
    wire _706 = 1'b0;
    wire _704 = 1'b0;
    wire _703 = 1'b0;
    wire _701 = 1'b0;
    wire _700 = 1'b0;
    wire _698 = 1'b0;
    wire _697 = 1'b0;
    wire _695 = 1'b0;
    wire _694 = 1'b0;
    reg _696;
    reg _699;
    reg _702;
    reg _705;
    reg _708;
    reg _711;
    reg _714;
    reg _717;
    reg _720;
    wire _749;
    wire _750;
    wire write_enable_34;
    wire _755;
    wire [131:0] _762;
    wire [63:0] _763;
    wire _691 = 1'b0;
    wire _690 = 1'b0;
    wire _693;
    wire _23;
    reg PHASE_7;
    wire [63:0] _775;
    wire [11:0] address_35;
    wire write_enable_35;
    wire [11:0] address_36;
    wire _962;
    wire read_enable_29;
    wire _960;
    wire write_enable_36;
    wire _964;
    wire [131:0] _969;
    wire [63:0] _970;
    wire [11:0] _955 = 12'b000000000000;
    wire [11:0] address_37;
    wire _953;
    wire write_enable_37;
    wire [63:0] _878;
    wire [63:0] _877;
    wire [63:0] _879;
    wire [63:0] _875;
    wire [63:0] _874;
    wire [63:0] q1_2;
    wire [63:0] _880;
    wire [11:0] address_38;
    wire write_enable_38 = 1'b0;
    wire _865;
    wire read_enable_30;
    wire [11:0] address_39;
    wire _861;
    wire read_enable_31;
    wire _859;
    wire write_enable_39;
    wire _863;
    wire [131:0] _870;
    wire [63:0] _871;
    wire [63:0] data_35 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_36;
    wire [11:0] _853 = 12'b000000000000;
    wire _851;
    wire _850;
    wire _849;
    wire _848;
    wire _847;
    wire _846;
    wire _845;
    wire _844;
    wire _843;
    wire _842;
    wire _841;
    wire _840;
    wire [11:0] _852;
    wire [11:0] address_40;
    wire write_enable_40 = 1'b0;
    wire _837;
    wire read_enable_32;
    wire [63:0] data_37;
    wire [63:0] data_38;
    wire _834;
    wire _833;
    wire _832;
    wire _831;
    wire _830;
    wire _829;
    wire _828;
    wire _827;
    wire _826;
    wire _825;
    wire _824;
    wire _823;
    wire [11:0] _835;
    wire [11:0] address_41;
    wire _820;
    wire read_enable_33;
    wire _818;
    wire write_enable_41;
    wire _822;
    wire [131:0] _857;
    wire [63:0] _858;
    wire _777 = 1'b0;
    wire _776 = 1'b0;
    wire _779;
    wire _27;
    reg PHASE_8;
    wire [63:0] _872;
    wire [11:0] address_42;
    wire _810;
    wire read_enable_34;
    wire write_enable_42;
    wire _812;
    wire [11:0] address_43;
    wire _805;
    wire read_enable_35;
    wire _803;
    wire write_enable_43;
    wire _807;
    wire [131:0] _815;
    wire [63:0] _816;
    wire [63:0] _883;
    wire [63:0] data_39;
    wire [63:0] data_40;
    wire [63:0] data_41;
    wire [63:0] data_42;
    wire [11:0] address_44;
    wire _796;
    wire read_enable_36;
    wire _793;
    wire _794;
    wire write_enable_44;
    wire _798;
    wire [11:0] address_45;
    wire _789;
    wire read_enable_37;
    wire _786;
    wire _787;
    wire write_enable_45;
    wire _791;
    wire [131:0] _801;
    wire [63:0] _802;
    wire _784 = 1'b0;
    wire _783 = 1'b0;
    wire _884;
    wire _29;
    reg PHASE_9;
    wire [63:0] q0_2;
    wire _781 = 1'b0;
    wire _780 = 1'b0;
    reg _782;
    wire [63:0] _873;
    wire [191:0] _882;
    wire [63:0] _885;
    wire [63:0] data_43;
    wire [63:0] data_44;
    wire [63:0] data_45;
    wire [63:0] data_46;
    wire [11:0] address_46;
    wire _949;
    wire _948;
    wire read_enable_38;
    wire _942 = 1'b0;
    wire _941 = 1'b0;
    wire _939 = 1'b0;
    wire _938 = 1'b0;
    wire _936 = 1'b0;
    wire _935 = 1'b0;
    wire _933 = 1'b0;
    wire _932 = 1'b0;
    wire _930 = 1'b0;
    wire _929 = 1'b0;
    wire _927 = 1'b0;
    wire _926 = 1'b0;
    wire _924 = 1'b0;
    wire _923 = 1'b0;
    wire _921 = 1'b0;
    wire _920 = 1'b0;
    wire _918 = 1'b0;
    wire _917 = 1'b0;
    reg _919;
    reg _922;
    reg _925;
    reg _928;
    reg _931;
    reg _934;
    reg _937;
    reg _940;
    reg _943;
    wire _944;
    wire _915 = 1'b0;
    wire _914 = 1'b0;
    wire _912 = 1'b0;
    wire _911 = 1'b0;
    wire _909 = 1'b0;
    wire _908 = 1'b0;
    wire _906 = 1'b0;
    wire _905 = 1'b0;
    wire _903 = 1'b0;
    wire _902 = 1'b0;
    wire _900 = 1'b0;
    wire _899 = 1'b0;
    wire _897 = 1'b0;
    wire _896 = 1'b0;
    wire _894 = 1'b0;
    wire _893 = 1'b0;
    wire _891 = 1'b0;
    wire _890 = 1'b0;
    reg _892;
    reg _895;
    reg _898;
    reg _901;
    reg _904;
    reg _907;
    reg _910;
    reg _913;
    reg _916;
    wire _945;
    wire _946;
    wire write_enable_46;
    wire _951;
    wire [131:0] _958;
    wire [63:0] _959;
    wire _887 = 1'b0;
    wire _886 = 1'b0;
    wire _889;
    wire _31;
    reg PHASE_10;
    wire [63:0] _971;
    wire [11:0] address_47;
    wire write_enable_47;
    wire [11:0] address_48;
    wire _1158;
    wire read_enable_39;
    wire _1156;
    wire write_enable_48;
    wire _1160;
    wire [131:0] _1165;
    wire [63:0] _1166;
    wire [11:0] _1151 = 12'b000000000000;
    wire [11:0] address_49;
    wire _1149;
    wire write_enable_49;
    wire [63:0] _1074;
    wire [63:0] _1073;
    wire [63:0] _1075;
    wire [63:0] _1071;
    wire [63:0] _1070;
    wire [63:0] q1_3;
    wire [63:0] _1076;
    wire [11:0] address_50;
    wire write_enable_50 = 1'b0;
    wire _1061;
    wire read_enable_40;
    wire [11:0] address_51;
    wire _1057;
    wire read_enable_41;
    wire _1055;
    wire write_enable_51;
    wire _1059;
    wire [131:0] _1066;
    wire [63:0] _1067;
    wire [63:0] data_47 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_48;
    wire [11:0] _1049 = 12'b000000000000;
    wire _1047;
    wire _1046;
    wire _1045;
    wire _1044;
    wire _1043;
    wire _1042;
    wire _1041;
    wire _1040;
    wire _1039;
    wire _1038;
    wire _1037;
    wire _1036;
    wire [11:0] _1048;
    wire [11:0] address_52;
    wire write_enable_52 = 1'b0;
    wire _1033;
    wire read_enable_42;
    wire [63:0] data_49;
    wire [63:0] data_50;
    wire _1030;
    wire _1029;
    wire _1028;
    wire _1027;
    wire _1026;
    wire _1025;
    wire _1024;
    wire _1023;
    wire _1022;
    wire _1021;
    wire _1020;
    wire _1019;
    wire [11:0] _1031;
    wire [11:0] address_53;
    wire _1016;
    wire read_enable_43;
    wire _1014;
    wire write_enable_53;
    wire _1018;
    wire [131:0] _1053;
    wire [63:0] _1054;
    wire _973 = 1'b0;
    wire _972 = 1'b0;
    wire _975;
    wire _35;
    reg PHASE_11;
    wire [63:0] _1068;
    wire [11:0] address_54;
    wire _1006;
    wire read_enable_44;
    wire write_enable_54;
    wire _1008;
    wire [11:0] address_55;
    wire _1001;
    wire read_enable_45;
    wire _999;
    wire write_enable_55;
    wire _1003;
    wire [131:0] _1011;
    wire [63:0] _1012;
    wire [63:0] _1079;
    wire [63:0] data_51;
    wire [63:0] data_52;
    wire [63:0] data_53;
    wire [63:0] data_54;
    wire [11:0] address_56;
    wire _992;
    wire read_enable_46;
    wire _989;
    wire _990;
    wire write_enable_56;
    wire _994;
    wire [11:0] address_57;
    wire _985;
    wire read_enable_47;
    wire _982;
    wire _983;
    wire write_enable_57;
    wire _987;
    wire [131:0] _997;
    wire [63:0] _998;
    wire _980 = 1'b0;
    wire _979 = 1'b0;
    wire _1080;
    wire _37;
    reg PHASE_12;
    wire [63:0] q0_3;
    wire _977 = 1'b0;
    wire _976 = 1'b0;
    reg _978;
    wire [63:0] _1069;
    wire [191:0] _1078;
    wire [63:0] _1081;
    wire [63:0] data_55;
    wire [63:0] data_56;
    wire [63:0] data_57;
    wire [63:0] data_58;
    wire [11:0] address_58;
    wire _1145;
    wire _1144;
    wire read_enable_48;
    wire _1138 = 1'b0;
    wire _1137 = 1'b0;
    wire _1135 = 1'b0;
    wire _1134 = 1'b0;
    wire _1132 = 1'b0;
    wire _1131 = 1'b0;
    wire _1129 = 1'b0;
    wire _1128 = 1'b0;
    wire _1126 = 1'b0;
    wire _1125 = 1'b0;
    wire _1123 = 1'b0;
    wire _1122 = 1'b0;
    wire _1120 = 1'b0;
    wire _1119 = 1'b0;
    wire _1117 = 1'b0;
    wire _1116 = 1'b0;
    wire _1114 = 1'b0;
    wire _1113 = 1'b0;
    reg _1115;
    reg _1118;
    reg _1121;
    reg _1124;
    reg _1127;
    reg _1130;
    reg _1133;
    reg _1136;
    reg _1139;
    wire _1140;
    wire _1111 = 1'b0;
    wire _1110 = 1'b0;
    wire _1108 = 1'b0;
    wire _1107 = 1'b0;
    wire _1105 = 1'b0;
    wire _1104 = 1'b0;
    wire _1102 = 1'b0;
    wire _1101 = 1'b0;
    wire _1099 = 1'b0;
    wire _1098 = 1'b0;
    wire _1096 = 1'b0;
    wire _1095 = 1'b0;
    wire _1093 = 1'b0;
    wire _1092 = 1'b0;
    wire _1090 = 1'b0;
    wire _1089 = 1'b0;
    wire _1087 = 1'b0;
    wire _1086 = 1'b0;
    reg _1088;
    reg _1091;
    reg _1094;
    reg _1097;
    reg _1100;
    reg _1103;
    reg _1106;
    reg _1109;
    reg _1112;
    wire _1141;
    wire _1142;
    wire write_enable_58;
    wire _1147;
    wire [131:0] _1154;
    wire [63:0] _1155;
    wire _1083 = 1'b0;
    wire _1082 = 1'b0;
    wire _1085;
    wire _39;
    reg PHASE_13;
    wire [63:0] _1167;
    wire [11:0] address_59;
    wire write_enable_59;
    wire [11:0] address_60;
    wire _1354;
    wire read_enable_49;
    wire _1352;
    wire write_enable_60;
    wire _1356;
    wire [131:0] _1361;
    wire [63:0] _1362;
    wire [11:0] _1347 = 12'b000000000000;
    wire [11:0] address_61;
    wire _1345;
    wire write_enable_61;
    wire [63:0] _1270;
    wire [63:0] _1269;
    wire [63:0] _1271;
    wire [63:0] _1267;
    wire [63:0] _1266;
    wire [63:0] q1_4;
    wire [63:0] _1272;
    wire [11:0] address_62;
    wire write_enable_62 = 1'b0;
    wire _1257;
    wire read_enable_50;
    wire [11:0] address_63;
    wire _1253;
    wire read_enable_51;
    wire _1251;
    wire write_enable_63;
    wire _1255;
    wire [131:0] _1262;
    wire [63:0] _1263;
    wire [63:0] data_59 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_60;
    wire [11:0] _1245 = 12'b000000000000;
    wire _1243;
    wire _1242;
    wire _1241;
    wire _1240;
    wire _1239;
    wire _1238;
    wire _1237;
    wire _1236;
    wire _1235;
    wire _1234;
    wire _1233;
    wire _1232;
    wire [11:0] _1244;
    wire [11:0] address_64;
    wire write_enable_64 = 1'b0;
    wire _1229;
    wire read_enable_52;
    wire [63:0] data_61;
    wire [63:0] data_62;
    wire _1226;
    wire _1225;
    wire _1224;
    wire _1223;
    wire _1222;
    wire _1221;
    wire _1220;
    wire _1219;
    wire _1218;
    wire _1217;
    wire _1216;
    wire _1215;
    wire [11:0] _1227;
    wire [11:0] address_65;
    wire _1212;
    wire read_enable_53;
    wire _1210;
    wire write_enable_65;
    wire _1214;
    wire [131:0] _1249;
    wire [63:0] _1250;
    wire _1169 = 1'b0;
    wire _1168 = 1'b0;
    wire _1171;
    wire _43;
    reg PHASE_14;
    wire [63:0] _1264;
    wire [11:0] address_66;
    wire _1202;
    wire read_enable_54;
    wire write_enable_66;
    wire _1204;
    wire [11:0] address_67;
    wire _1197;
    wire read_enable_55;
    wire _1195;
    wire write_enable_67;
    wire _1199;
    wire [131:0] _1207;
    wire [63:0] _1208;
    wire [63:0] _1275;
    wire [63:0] data_63;
    wire [63:0] data_64;
    wire [63:0] data_65;
    wire [63:0] data_66;
    wire [11:0] address_68;
    wire _1188;
    wire read_enable_56;
    wire _1185;
    wire _1186;
    wire write_enable_68;
    wire _1190;
    wire [11:0] address_69;
    wire _1181;
    wire read_enable_57;
    wire _1178;
    wire _1179;
    wire write_enable_69;
    wire _1183;
    wire [131:0] _1193;
    wire [63:0] _1194;
    wire _1176 = 1'b0;
    wire _1175 = 1'b0;
    wire _1276;
    wire _45;
    reg PHASE_15;
    wire [63:0] q0_4;
    wire _1173 = 1'b0;
    wire _1172 = 1'b0;
    reg _1174;
    wire [63:0] _1265;
    wire [191:0] _1274;
    wire [63:0] _1277;
    wire [63:0] data_67;
    wire [63:0] data_68;
    wire [63:0] data_69;
    wire [63:0] data_70;
    wire [11:0] address_70;
    wire _1341;
    wire _1340;
    wire read_enable_58;
    wire _1334 = 1'b0;
    wire _1333 = 1'b0;
    wire _1331 = 1'b0;
    wire _1330 = 1'b0;
    wire _1328 = 1'b0;
    wire _1327 = 1'b0;
    wire _1325 = 1'b0;
    wire _1324 = 1'b0;
    wire _1322 = 1'b0;
    wire _1321 = 1'b0;
    wire _1319 = 1'b0;
    wire _1318 = 1'b0;
    wire _1316 = 1'b0;
    wire _1315 = 1'b0;
    wire _1313 = 1'b0;
    wire _1312 = 1'b0;
    wire _1310 = 1'b0;
    wire _1309 = 1'b0;
    reg _1311;
    reg _1314;
    reg _1317;
    reg _1320;
    reg _1323;
    reg _1326;
    reg _1329;
    reg _1332;
    reg _1335;
    wire _1336;
    wire _1307 = 1'b0;
    wire _1306 = 1'b0;
    wire _1304 = 1'b0;
    wire _1303 = 1'b0;
    wire _1301 = 1'b0;
    wire _1300 = 1'b0;
    wire _1298 = 1'b0;
    wire _1297 = 1'b0;
    wire _1295 = 1'b0;
    wire _1294 = 1'b0;
    wire _1292 = 1'b0;
    wire _1291 = 1'b0;
    wire _1289 = 1'b0;
    wire _1288 = 1'b0;
    wire _1286 = 1'b0;
    wire _1285 = 1'b0;
    wire _1283 = 1'b0;
    wire _1282 = 1'b0;
    reg _1284;
    reg _1287;
    reg _1290;
    reg _1293;
    reg _1296;
    reg _1299;
    reg _1302;
    reg _1305;
    reg _1308;
    wire _1337;
    wire _1338;
    wire write_enable_70;
    wire _1343;
    wire [131:0] _1350;
    wire [63:0] _1351;
    wire _1279 = 1'b0;
    wire _1278 = 1'b0;
    wire _1281;
    wire _47;
    reg PHASE_16;
    wire [63:0] _1363;
    wire [11:0] address_71;
    wire write_enable_71;
    wire [11:0] address_72;
    wire _1550;
    wire read_enable_59;
    wire _1548;
    wire write_enable_72;
    wire _1552;
    wire [131:0] _1557;
    wire [63:0] _1558;
    wire [11:0] _1543 = 12'b000000000000;
    wire [11:0] address_73;
    wire _1541;
    wire write_enable_73;
    wire [63:0] _1466;
    wire [63:0] _1465;
    wire [63:0] _1467;
    wire [63:0] _1463;
    wire [63:0] _1462;
    wire [63:0] q1_5;
    wire [63:0] _1468;
    wire [11:0] address_74;
    wire write_enable_74 = 1'b0;
    wire _1453;
    wire read_enable_60;
    wire [11:0] address_75;
    wire _1449;
    wire read_enable_61;
    wire _1447;
    wire write_enable_75;
    wire _1451;
    wire [131:0] _1458;
    wire [63:0] _1459;
    wire [63:0] data_71 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_72;
    wire [11:0] _1441 = 12'b000000000000;
    wire _1439;
    wire _1438;
    wire _1437;
    wire _1436;
    wire _1435;
    wire _1434;
    wire _1433;
    wire _1432;
    wire _1431;
    wire _1430;
    wire _1429;
    wire _1428;
    wire [11:0] _1440;
    wire [11:0] address_76;
    wire write_enable_76 = 1'b0;
    wire _1425;
    wire read_enable_62;
    wire [63:0] data_73;
    wire [63:0] data_74;
    wire _1422;
    wire _1421;
    wire _1420;
    wire _1419;
    wire _1418;
    wire _1417;
    wire _1416;
    wire _1415;
    wire _1414;
    wire _1413;
    wire _1412;
    wire _1411;
    wire [11:0] _1423;
    wire [11:0] address_77;
    wire _1408;
    wire read_enable_63;
    wire _1406;
    wire write_enable_77;
    wire _1410;
    wire [131:0] _1445;
    wire [63:0] _1446;
    wire _1365 = 1'b0;
    wire _1364 = 1'b0;
    wire _1367;
    wire _51;
    reg PHASE_17;
    wire [63:0] _1460;
    wire [11:0] address_78;
    wire _1398;
    wire read_enable_64;
    wire write_enable_78;
    wire _1400;
    wire [11:0] address_79;
    wire _1393;
    wire read_enable_65;
    wire _1391;
    wire write_enable_79;
    wire _1395;
    wire [131:0] _1403;
    wire [63:0] _1404;
    wire [63:0] _1471;
    wire [63:0] data_75;
    wire [63:0] data_76;
    wire [63:0] data_77;
    wire [63:0] data_78;
    wire [11:0] address_80;
    wire _1384;
    wire read_enable_66;
    wire _1381;
    wire _1382;
    wire write_enable_80;
    wire _1386;
    wire [11:0] address_81;
    wire _1377;
    wire read_enable_67;
    wire _1374;
    wire _1375;
    wire write_enable_81;
    wire _1379;
    wire [131:0] _1389;
    wire [63:0] _1390;
    wire _1372 = 1'b0;
    wire _1371 = 1'b0;
    wire _1472;
    wire _53;
    reg PHASE_18;
    wire [63:0] q0_5;
    wire _1369 = 1'b0;
    wire _1368 = 1'b0;
    reg _1370;
    wire [63:0] _1461;
    wire [191:0] _1470;
    wire [63:0] _1473;
    wire [63:0] data_79;
    wire [63:0] data_80;
    wire [63:0] data_81;
    wire [63:0] data_82;
    wire [11:0] address_82;
    wire _1537;
    wire _1536;
    wire read_enable_68;
    wire _1530 = 1'b0;
    wire _1529 = 1'b0;
    wire _1527 = 1'b0;
    wire _1526 = 1'b0;
    wire _1524 = 1'b0;
    wire _1523 = 1'b0;
    wire _1521 = 1'b0;
    wire _1520 = 1'b0;
    wire _1518 = 1'b0;
    wire _1517 = 1'b0;
    wire _1515 = 1'b0;
    wire _1514 = 1'b0;
    wire _1512 = 1'b0;
    wire _1511 = 1'b0;
    wire _1509 = 1'b0;
    wire _1508 = 1'b0;
    wire _1506 = 1'b0;
    wire _1505 = 1'b0;
    reg _1507;
    reg _1510;
    reg _1513;
    reg _1516;
    reg _1519;
    reg _1522;
    reg _1525;
    reg _1528;
    reg _1531;
    wire _1532;
    wire _1503 = 1'b0;
    wire _1502 = 1'b0;
    wire _1500 = 1'b0;
    wire _1499 = 1'b0;
    wire _1497 = 1'b0;
    wire _1496 = 1'b0;
    wire _1494 = 1'b0;
    wire _1493 = 1'b0;
    wire _1491 = 1'b0;
    wire _1490 = 1'b0;
    wire _1488 = 1'b0;
    wire _1487 = 1'b0;
    wire _1485 = 1'b0;
    wire _1484 = 1'b0;
    wire _1482 = 1'b0;
    wire _1481 = 1'b0;
    wire _1479 = 1'b0;
    wire _1478 = 1'b0;
    reg _1480;
    reg _1483;
    reg _1486;
    reg _1489;
    reg _1492;
    reg _1495;
    reg _1498;
    reg _1501;
    reg _1504;
    wire _1533;
    wire _1534;
    wire write_enable_82;
    wire _1539;
    wire [131:0] _1546;
    wire [63:0] _1547;
    wire _1475 = 1'b0;
    wire _1474 = 1'b0;
    wire _1477;
    wire _55;
    reg PHASE_19;
    wire [63:0] _1559;
    wire [11:0] address_83;
    wire write_enable_83;
    wire [11:0] address_84;
    wire _1746;
    wire read_enable_69;
    wire _1744;
    wire write_enable_84;
    wire _1748;
    wire [131:0] _1753;
    wire [63:0] _1754;
    wire [11:0] _1739 = 12'b000000000000;
    wire [11:0] address_85;
    wire _1737;
    wire write_enable_85;
    wire [3:0] _292;
    wire _291;
    wire _289;
    wire [63:0] _288;
    wire [63:0] _287;
    wire [63:0] _286;
    wire [63:0] _285;
    wire [63:0] _284;
    wire [63:0] _283;
    wire [63:0] _282;
    wire [63:0] _1662;
    wire [63:0] _1661;
    wire [63:0] _1663;
    wire [63:0] _1659;
    wire [63:0] _1658;
    wire [63:0] q1_6;
    wire [63:0] _1664;
    wire [11:0] address_86;
    wire write_enable_86 = 1'b0;
    wire _1649;
    wire read_enable_70;
    wire [11:0] address_87;
    wire _1645;
    wire read_enable_71;
    wire _1643;
    wire write_enable_87;
    wire _1647;
    wire [131:0] _1654;
    wire [63:0] _1655;
    wire [63:0] data_83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_84;
    wire [11:0] _1637 = 12'b000000000000;
    wire _1635;
    wire _1634;
    wire _1633;
    wire _1632;
    wire _1631;
    wire _1630;
    wire _1629;
    wire _1628;
    wire _1627;
    wire _1626;
    wire _1625;
    wire _1624;
    wire [11:0] _1636;
    wire [11:0] address_88;
    wire write_enable_88 = 1'b0;
    wire _1621;
    wire read_enable_72;
    wire [63:0] data_85;
    wire [63:0] data_86;
    wire [11:0] _60;
    wire _1618;
    wire _1617;
    wire _1616;
    wire _1615;
    wire _1614;
    wire _1613;
    wire _1612;
    wire _1611;
    wire _1610;
    wire _1609;
    wire _1608;
    wire _1607;
    wire [11:0] _1619;
    wire [11:0] address_89;
    wire _1604;
    wire read_enable_73;
    wire [7:0] _62;
    wire _1602;
    wire write_enable_89;
    wire _1606;
    wire [131:0] _1641;
    wire [63:0] _1642;
    wire _1561 = 1'b0;
    wire _1560 = 1'b0;
    wire _1563;
    wire _63;
    reg PHASE_20;
    wire [63:0] _1656;
    wire [11:0] address_90;
    wire _1594;
    wire read_enable_74;
    wire write_enable_90;
    wire _1596;
    wire [11:0] address_91;
    wire _1589;
    wire read_enable_75;
    wire _1587;
    wire write_enable_91;
    wire _1591;
    wire [131:0] _1599;
    wire [63:0] _1600;
    wire [63:0] _1667;
    wire [63:0] data_87;
    wire [63:0] data_88;
    wire [63:0] data_89;
    wire [63:0] data_90;
    wire [11:0] _198 = 12'b000000000000;
    wire [11:0] _197 = 12'b000000000000;
    wire [11:0] _195 = 12'b000000000000;
    wire [11:0] _194 = 12'b000000000000;
    wire [11:0] _192 = 12'b000000000000;
    wire [11:0] _191 = 12'b000000000000;
    wire [11:0] _189 = 12'b000000000000;
    wire [11:0] _188 = 12'b000000000000;
    wire [11:0] _186 = 12'b000000000000;
    wire [11:0] _185 = 12'b000000000000;
    wire [11:0] _183 = 12'b000000000000;
    wire [11:0] _182 = 12'b000000000000;
    wire [11:0] _180 = 12'b000000000000;
    wire [11:0] _179 = 12'b000000000000;
    wire [11:0] _177 = 12'b000000000000;
    wire [11:0] _176 = 12'b000000000000;
    wire [11:0] _174 = 12'b000000000000;
    wire [11:0] _173 = 12'b000000000000;
    reg [11:0] _175;
    reg [11:0] _178;
    reg [11:0] _181;
    reg [11:0] _184;
    reg [11:0] _187;
    reg [11:0] _190;
    reg [11:0] _193;
    reg [11:0] _196;
    reg [11:0] _199;
    wire [11:0] _172;
    wire [11:0] address_92;
    wire _1580;
    wire read_enable_76;
    wire _1577;
    wire _1578;
    wire write_enable_92;
    wire _1582;
    wire [11:0] address_93;
    wire _1573;
    wire read_enable_77;
    wire _1570;
    wire _1571;
    wire write_enable_93;
    wire _1575;
    wire [131:0] _1585;
    wire [63:0] _1586;
    wire _99;
    wire _1568 = 1'b0;
    wire _1567 = 1'b0;
    wire _1668;
    wire _65;
    reg PHASE_21;
    wire [63:0] q0_6;
    wire _1565 = 1'b0;
    wire _1564 = 1'b0;
    wire _92;
    reg _1566;
    wire [63:0] _1657;
    wire [191:0] _1666;
    wire [63:0] _1669;
    wire [63:0] data_91;
    wire [63:0] data_92;
    wire [63:0] data_93;
    wire [63:0] data_94;
    wire [11:0] _163 = 12'b000000000000;
    wire [11:0] _162 = 12'b000000000000;
    wire [11:0] _160 = 12'b000000000000;
    wire [11:0] _159 = 12'b000000000000;
    wire [11:0] _157 = 12'b000000000000;
    wire [11:0] _156 = 12'b000000000000;
    wire [11:0] _154 = 12'b000000000000;
    wire [11:0] _153 = 12'b000000000000;
    wire [11:0] _151 = 12'b000000000000;
    wire [11:0] _150 = 12'b000000000000;
    wire [11:0] _148 = 12'b000000000000;
    wire [11:0] _147 = 12'b000000000000;
    wire [11:0] _145 = 12'b000000000000;
    wire [11:0] _144 = 12'b000000000000;
    wire [11:0] _142 = 12'b000000000000;
    wire [11:0] _141 = 12'b000000000000;
    wire [11:0] _139 = 12'b000000000000;
    wire [11:0] _138 = 12'b000000000000;
    wire [11:0] _137;
    reg [11:0] _140;
    reg [11:0] _143;
    reg [11:0] _146;
    reg [11:0] _149;
    reg [11:0] _152;
    reg [11:0] _155;
    reg [11:0] _158;
    reg [11:0] _161;
    reg [11:0] _164;
    wire [11:0] _68;
    wire [11:0] address_94;
    wire _1733;
    wire [7:0] _70;
    wire _1732;
    wire read_enable_78;
    wire _1726 = 1'b0;
    wire _1725 = 1'b0;
    wire _1723 = 1'b0;
    wire _1722 = 1'b0;
    wire _1720 = 1'b0;
    wire _1719 = 1'b0;
    wire _1717 = 1'b0;
    wire _1716 = 1'b0;
    wire _1714 = 1'b0;
    wire _1713 = 1'b0;
    wire _1711 = 1'b0;
    wire _1710 = 1'b0;
    wire _1708 = 1'b0;
    wire _1707 = 1'b0;
    wire _1705 = 1'b0;
    wire _1704 = 1'b0;
    wire _1702 = 1'b0;
    wire _1701 = 1'b0;
    wire _290;
    reg _1703;
    reg _1706;
    reg _1709;
    reg _1712;
    reg _1715;
    reg _1718;
    reg _1721;
    reg _1724;
    reg _1727;
    wire _1728;
    wire _1699 = 1'b0;
    wire _1698 = 1'b0;
    wire _1696 = 1'b0;
    wire _1695 = 1'b0;
    wire _1693 = 1'b0;
    wire _1692 = 1'b0;
    wire _1690 = 1'b0;
    wire _1689 = 1'b0;
    wire _1687 = 1'b0;
    wire _1686 = 1'b0;
    wire _1684 = 1'b0;
    wire _1683 = 1'b0;
    wire _1681 = 1'b0;
    wire _1680 = 1'b0;
    wire _1678 = 1'b0;
    wire _1677 = 1'b0;
    wire _1675 = 1'b0;
    wire _1674 = 1'b0;
    wire _130;
    reg _1676;
    reg _1679;
    reg _1682;
    reg _1685;
    reg _1688;
    reg _1691;
    reg _1694;
    reg _1697;
    reg _1700;
    wire _1729;
    wire _128 = 1'b0;
    wire _127 = 1'b0;
    wire _125 = 1'b0;
    wire _124 = 1'b0;
    wire _122 = 1'b0;
    wire _121 = 1'b0;
    wire _119 = 1'b0;
    wire _118 = 1'b0;
    wire _116 = 1'b0;
    wire _115 = 1'b0;
    wire _113 = 1'b0;
    wire _112 = 1'b0;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire vdd = 1'b1;
    wire _104 = 1'b0;
    wire _103 = 1'b0;
    wire _102;
    reg _105;
    reg _108;
    reg _111;
    reg _114;
    reg _117;
    reg _120;
    reg _123;
    reg _126;
    reg _129;
    wire _1730;
    wire write_enable_94;
    wire _1735;
    wire gnd = 1'b0;
    wire [131:0] _1742;
    wire [63:0] _1743;
    wire _72;
    wire _1671 = 1'b0;
    wire _1670 = 1'b0;
    wire _1673;
    wire _73;
    reg PHASE_22;
    wire [63:0] _1755;
    wire _76;
    wire _78;
    wire _80;
    wire _82;
    wire _84;
    wire [523:0] _91;
    wire _1756;

    /* logic */
    assign address = _372 ? _199 : _367;
    assign write_enable = _365 & _372;
    assign address_0 = _372 ? _164 : _68;
    assign _374 = ~ _372;
    assign read_enable = _360 & _374;
    assign _372 = ~ PHASE_1;
    assign write_enable_0 = _358 & _372;
    assign _376 = write_enable_0 | read_enable;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_376), .regcea(vdd), .wea(write_enable_0), .addra(address_0), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable), .regceb(vdd), .web(write_enable), .addrb(address), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_381[131:131]), .sbiterrb(_381[130:130]), .doutb(_381[129:66]), .dbiterra(_381[65:65]), .sbiterra(_381[64:64]), .douta(_381[63:0]) );
    assign _382 = _381[63:0];
    assign address_1 = PHASE_1 ? _199 : _367;
    assign _365 = _129 & _328;
    assign write_enable_1 = _365 & PHASE_1;
    assign _279 = _271[129:66];
    assign _278 = _258[129:66];
    assign _280 = PHASE ? _279 : _278;
    assign _276 = _216[129:66];
    assign _275 = _202[129:66];
    assign q1 = PHASE_0 ? _276 : _275;
    assign _281 = _96 ? _280 : q1;
    assign address_2 = _260 ? _254 : _253;
    assign _266 = ~ _260;
    assign read_enable_0 = _102 & _266;
    assign address_3 = _260 ? _60 : _236;
    assign _262 = ~ _260;
    assign read_enable_1 = _102 & _262;
    assign _260 = ~ PHASE;
    assign write_enable_3 = _219 & _260;
    assign _264 = write_enable_3 | read_enable_1;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_0
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_264), .regcea(vdd), .wea(write_enable_3), .addra(address_3), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_0), .regceb(vdd), .web(write_enable_2), .addrb(address_2), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_271[131:131]), .sbiterrb(_271[130:130]), .doutb(_271[129:66]), .dbiterra(_271[65:65]), .sbiterra(_271[64:64]), .douta(_271[63:0]) );
    assign _272 = _271[63:0];
    assign _252 = _172[11:11];
    assign _251 = _172[10:10];
    assign _250 = _172[9:9];
    assign _249 = _172[8:8];
    assign _248 = _172[7:7];
    assign _247 = _172[6:6];
    assign _246 = _172[5:5];
    assign _245 = _172[4:4];
    assign _244 = _172[3:3];
    assign _243 = _172[2:2];
    assign _242 = _172[1:1];
    assign _241 = _172[0:0];
    assign _253 = { _241, _242, _243, _244, _245, _246, _247, _248, _249, _250, _251, _252 };
    assign address_4 = PHASE ? _254 : _253;
    assign _238 = ~ PHASE;
    assign read_enable_2 = _102 & _238;
    assign data_1 = wr_d7;
    assign _235 = _137[11:11];
    assign _234 = _137[10:10];
    assign _233 = _137[9:9];
    assign _232 = _137[8:8];
    assign _231 = _137[7:7];
    assign _230 = _137[6:6];
    assign _229 = _137[5:5];
    assign _228 = _137[4:4];
    assign _227 = _137[3:3];
    assign _226 = _137[2:2];
    assign _225 = _137[1:1];
    assign _224 = _137[0:0];
    assign _236 = { _224, _225, _226, _227, _228, _229, _230, _231, _232, _233, _234, _235 };
    assign address_5 = PHASE ? _60 : _236;
    assign _221 = ~ PHASE;
    assign read_enable_3 = _102 & _221;
    assign _219 = _62[7:7];
    assign write_enable_5 = _219 & PHASE;
    assign _223 = write_enable_5 | read_enable_3;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_1
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_223), .regcea(vdd), .wea(write_enable_5), .addra(address_5), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_2), .regceb(vdd), .web(write_enable_4), .addrb(address_4), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_258[131:131]), .sbiterrb(_258[130:130]), .doutb(_258[129:66]), .dbiterra(_258[65:65]), .sbiterra(_258[64:64]), .douta(_258[63:0]) );
    assign _259 = _258[63:0];
    assign _89 = ~ PHASE;
    assign _3 = _89;
    always @(posedge _84) begin
        if (_82)
            PHASE <= _87;
        else
            if (_72)
                PHASE <= _3;
    end
    assign _273 = PHASE ? _272 : _259;
    assign address_6 = _204 ? _199 : _172;
    assign _211 = ~ _204;
    assign read_enable_4 = _102 & _211;
    assign write_enable_6 = _167 & _204;
    assign _213 = write_enable_6 | read_enable_4;
    assign address_7 = _204 ? _164 : _137;
    assign _206 = ~ _204;
    assign read_enable_5 = _102 & _206;
    assign _204 = ~ PHASE_0;
    assign write_enable_7 = _132 & _204;
    assign _208 = write_enable_7 | read_enable_5;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_2
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_208), .regcea(vdd), .wea(write_enable_7), .addra(address_7), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_213), .regceb(vdd), .web(write_enable_6), .addrb(address_6), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_216[131:131]), .sbiterrb(_216[130:130]), .doutb(_216[129:66]), .dbiterra(_216[65:65]), .sbiterra(_216[64:64]), .douta(_216[63:0]) );
    assign _217 = _216[63:0];
    assign _295 = _294[127:64];
    assign data_3 = _295;
    assign address_8 = PHASE_0 ? _199 : _172;
    assign _169 = ~ PHASE_0;
    assign read_enable_6 = _102 & _169;
    assign _166 = ~ _130;
    assign _167 = _129 & _166;
    assign write_enable_8 = _167 & PHASE_0;
    assign _171 = write_enable_8 | read_enable_6;
    assign address_9 = PHASE_0 ? _164 : _137;
    assign _134 = ~ PHASE_0;
    assign read_enable_7 = _102 & _134;
    assign _131 = ~ _130;
    assign _132 = _129 & _131;
    assign write_enable_9 = _132 & PHASE_0;
    assign _136 = write_enable_9 | read_enable_7;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_3
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_136), .regcea(vdd), .wea(write_enable_9), .addra(address_9), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_171), .regceb(vdd), .web(write_enable_8), .addrb(address_8), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_202[131:131]), .sbiterrb(_202[130:130]), .doutb(_202[129:66]), .dbiterra(_202[65:65]), .sbiterra(_202[64:64]), .douta(_202[63:0]) );
    assign _203 = _202[63:0];
    assign _296 = ~ PHASE_0;
    assign _5 = _296;
    always @(posedge _84) begin
        if (_82)
            PHASE_0 <= _98;
        else
            if (_99)
                PHASE_0 <= _5;
    end
    assign q0 = PHASE_0 ? _217 : _203;
    always @(posedge _84) begin
        if (_82)
            _96 <= _94;
        else
            _96 <= _92;
    end
    assign _274 = _96 ? _273 : q0;
    dp_54
        dp_6
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_274), .d2(_281), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_294[191:128]), .q2(_294[127:64]), .q1(_294[63:0]) );
    assign _297 = _294[63:0];
    assign data_7 = _297;
    assign address_10 = PHASE_1 ? _164 : _68;
    assign _361 = ~ PHASE_1;
    assign _360 = _70[7:7];
    assign read_enable_8 = _360 & _361;
    always @(posedge _84) begin
        if (_82)
            _331 <= _330;
        else
            _331 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _334 <= _333;
        else
            _334 <= _331;
    end
    always @(posedge _84) begin
        if (_82)
            _337 <= _336;
        else
            _337 <= _334;
    end
    always @(posedge _84) begin
        if (_82)
            _340 <= _339;
        else
            _340 <= _337;
    end
    always @(posedge _84) begin
        if (_82)
            _343 <= _342;
        else
            _343 <= _340;
    end
    always @(posedge _84) begin
        if (_82)
            _346 <= _345;
        else
            _346 <= _343;
    end
    always @(posedge _84) begin
        if (_82)
            _349 <= _348;
        else
            _349 <= _346;
    end
    always @(posedge _84) begin
        if (_82)
            _352 <= _351;
        else
            _352 <= _349;
    end
    always @(posedge _84) begin
        if (_82)
            _355 <= _354;
        else
            _355 <= _352;
    end
    assign _356 = ~ _355;
    always @(posedge _84) begin
        if (_82)
            _304 <= _303;
        else
            _304 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _307 <= _306;
        else
            _307 <= _304;
    end
    always @(posedge _84) begin
        if (_82)
            _310 <= _309;
        else
            _310 <= _307;
    end
    always @(posedge _84) begin
        if (_82)
            _313 <= _312;
        else
            _313 <= _310;
    end
    always @(posedge _84) begin
        if (_82)
            _316 <= _315;
        else
            _316 <= _313;
    end
    always @(posedge _84) begin
        if (_82)
            _319 <= _318;
        else
            _319 <= _316;
    end
    always @(posedge _84) begin
        if (_82)
            _322 <= _321;
        else
            _322 <= _319;
    end
    always @(posedge _84) begin
        if (_82)
            _325 <= _324;
        else
            _325 <= _322;
    end
    always @(posedge _84) begin
        if (_82)
            _328 <= _327;
        else
            _328 <= _325;
    end
    assign _357 = _328 & _356;
    assign _358 = _129 & _357;
    assign write_enable_10 = _358 & PHASE_1;
    assign _363 = write_enable_10 | read_enable_8;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_4
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_363), .regcea(vdd), .wea(write_enable_10), .addra(address_10), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_1), .regceb(vdd), .web(write_enable_1), .addrb(address_1), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_370[131:131]), .sbiterrb(_370[130:130]), .doutb(_370[129:66]), .dbiterra(_370[65:65]), .sbiterra(_370[64:64]), .douta(_370[63:0]) );
    assign _371 = _370[63:0];
    assign _301 = ~ PHASE_1;
    assign _7 = _301;
    always @(posedge _84) begin
        if (_82)
            PHASE_1 <= _299;
        else
            if (_72)
                PHASE_1 <= _7;
    end
    assign _383 = PHASE_1 ? _382 : _371;
    assign address_11 = _568 ? _199 : _563;
    assign write_enable_11 = _561 & _568;
    assign address_12 = _568 ? _164 : _68;
    assign _570 = ~ _568;
    assign read_enable_9 = _556 & _570;
    assign _568 = ~ PHASE_4;
    assign write_enable_12 = _554 & _568;
    assign _572 = write_enable_12 | read_enable_9;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_5
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_572), .regcea(vdd), .wea(write_enable_12), .addra(address_12), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_11), .regceb(vdd), .web(write_enable_11), .addrb(address_11), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_577[131:131]), .sbiterrb(_577[130:130]), .doutb(_577[129:66]), .dbiterra(_577[65:65]), .sbiterra(_577[64:64]), .douta(_577[63:0]) );
    assign _578 = _577[63:0];
    assign address_13 = PHASE_4 ? _199 : _563;
    assign _561 = _129 & _524;
    assign write_enable_13 = _561 & PHASE_4;
    assign _486 = _478[129:66];
    assign _485 = _465[129:66];
    assign _487 = PHASE_2 ? _486 : _485;
    assign _483 = _423[129:66];
    assign _482 = _409[129:66];
    assign q1_0 = PHASE_3 ? _483 : _482;
    assign _488 = _390 ? _487 : q1_0;
    assign address_14 = _467 ? _461 : _460;
    assign _473 = ~ _467;
    assign read_enable_10 = _102 & _473;
    assign address_15 = _467 ? _60 : _443;
    assign _469 = ~ _467;
    assign read_enable_11 = _102 & _469;
    assign _467 = ~ PHASE_2;
    assign write_enable_15 = _426 & _467;
    assign _471 = write_enable_15 | read_enable_11;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_6
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_471), .regcea(vdd), .wea(write_enable_15), .addra(address_15), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_10), .regceb(vdd), .web(write_enable_14), .addrb(address_14), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_478[131:131]), .sbiterrb(_478[130:130]), .doutb(_478[129:66]), .dbiterra(_478[65:65]), .sbiterra(_478[64:64]), .douta(_478[63:0]) );
    assign _479 = _478[63:0];
    assign _459 = _172[11:11];
    assign _458 = _172[10:10];
    assign _457 = _172[9:9];
    assign _456 = _172[8:8];
    assign _455 = _172[7:7];
    assign _454 = _172[6:6];
    assign _453 = _172[5:5];
    assign _452 = _172[4:4];
    assign _451 = _172[3:3];
    assign _450 = _172[2:2];
    assign _449 = _172[1:1];
    assign _448 = _172[0:0];
    assign _460 = { _448, _449, _450, _451, _452, _453, _454, _455, _456, _457, _458, _459 };
    assign address_16 = PHASE_2 ? _461 : _460;
    assign _445 = ~ PHASE_2;
    assign read_enable_12 = _102 & _445;
    assign data_13 = wr_d6;
    assign _442 = _137[11:11];
    assign _441 = _137[10:10];
    assign _440 = _137[9:9];
    assign _439 = _137[8:8];
    assign _438 = _137[7:7];
    assign _437 = _137[6:6];
    assign _436 = _137[5:5];
    assign _435 = _137[4:4];
    assign _434 = _137[3:3];
    assign _433 = _137[2:2];
    assign _432 = _137[1:1];
    assign _431 = _137[0:0];
    assign _443 = { _431, _432, _433, _434, _435, _436, _437, _438, _439, _440, _441, _442 };
    assign address_17 = PHASE_2 ? _60 : _443;
    assign _428 = ~ PHASE_2;
    assign read_enable_13 = _102 & _428;
    assign _426 = _62[6:6];
    assign write_enable_17 = _426 & PHASE_2;
    assign _430 = write_enable_17 | read_enable_13;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_7
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_430), .regcea(vdd), .wea(write_enable_17), .addra(address_17), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_12), .regceb(vdd), .web(write_enable_16), .addrb(address_16), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_465[131:131]), .sbiterrb(_465[130:130]), .doutb(_465[129:66]), .dbiterra(_465[65:65]), .sbiterra(_465[64:64]), .douta(_465[63:0]) );
    assign _466 = _465[63:0];
    assign _387 = ~ PHASE_2;
    assign _11 = _387;
    always @(posedge _84) begin
        if (_82)
            PHASE_2 <= _385;
        else
            if (_72)
                PHASE_2 <= _11;
    end
    assign _480 = PHASE_2 ? _479 : _466;
    assign address_18 = _411 ? _199 : _172;
    assign _418 = ~ _411;
    assign read_enable_14 = _102 & _418;
    assign write_enable_18 = _402 & _411;
    assign _420 = write_enable_18 | read_enable_14;
    assign address_19 = _411 ? _164 : _137;
    assign _413 = ~ _411;
    assign read_enable_15 = _102 & _413;
    assign _411 = ~ PHASE_3;
    assign write_enable_19 = _395 & _411;
    assign _415 = write_enable_19 | read_enable_15;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_8
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_415), .regcea(vdd), .wea(write_enable_19), .addra(address_19), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_420), .regceb(vdd), .web(write_enable_18), .addrb(address_18), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_423[131:131]), .sbiterrb(_423[130:130]), .doutb(_423[129:66]), .dbiterra(_423[65:65]), .sbiterra(_423[64:64]), .douta(_423[63:0]) );
    assign _424 = _423[63:0];
    assign _491 = _490[127:64];
    assign data_15 = _491;
    assign address_20 = PHASE_3 ? _199 : _172;
    assign _404 = ~ PHASE_3;
    assign read_enable_16 = _102 & _404;
    assign _401 = ~ _130;
    assign _402 = _129 & _401;
    assign write_enable_20 = _402 & PHASE_3;
    assign _406 = write_enable_20 | read_enable_16;
    assign address_21 = PHASE_3 ? _164 : _137;
    assign _397 = ~ PHASE_3;
    assign read_enable_17 = _102 & _397;
    assign _394 = ~ _130;
    assign _395 = _129 & _394;
    assign write_enable_21 = _395 & PHASE_3;
    assign _399 = write_enable_21 | read_enable_17;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_9
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_399), .regcea(vdd), .wea(write_enable_21), .addra(address_21), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_406), .regceb(vdd), .web(write_enable_20), .addrb(address_20), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_409[131:131]), .sbiterrb(_409[130:130]), .doutb(_409[129:66]), .dbiterra(_409[65:65]), .sbiterra(_409[64:64]), .douta(_409[63:0]) );
    assign _410 = _409[63:0];
    assign _492 = ~ PHASE_3;
    assign _13 = _492;
    always @(posedge _84) begin
        if (_82)
            PHASE_3 <= _392;
        else
            if (_99)
                PHASE_3 <= _13;
    end
    assign q0_0 = PHASE_3 ? _424 : _410;
    always @(posedge _84) begin
        if (_82)
            _390 <= _389;
        else
            _390 <= _92;
    end
    assign _481 = _390 ? _480 : q0_0;
    dp_53
        dp_5
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_481), .d2(_488), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_490[191:128]), .q2(_490[127:64]), .q1(_490[63:0]) );
    assign _493 = _490[63:0];
    assign data_19 = _493;
    assign address_22 = PHASE_4 ? _164 : _68;
    assign _557 = ~ PHASE_4;
    assign _556 = _70[6:6];
    assign read_enable_18 = _556 & _557;
    always @(posedge _84) begin
        if (_82)
            _527 <= _526;
        else
            _527 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _530 <= _529;
        else
            _530 <= _527;
    end
    always @(posedge _84) begin
        if (_82)
            _533 <= _532;
        else
            _533 <= _530;
    end
    always @(posedge _84) begin
        if (_82)
            _536 <= _535;
        else
            _536 <= _533;
    end
    always @(posedge _84) begin
        if (_82)
            _539 <= _538;
        else
            _539 <= _536;
    end
    always @(posedge _84) begin
        if (_82)
            _542 <= _541;
        else
            _542 <= _539;
    end
    always @(posedge _84) begin
        if (_82)
            _545 <= _544;
        else
            _545 <= _542;
    end
    always @(posedge _84) begin
        if (_82)
            _548 <= _547;
        else
            _548 <= _545;
    end
    always @(posedge _84) begin
        if (_82)
            _551 <= _550;
        else
            _551 <= _548;
    end
    assign _552 = ~ _551;
    always @(posedge _84) begin
        if (_82)
            _500 <= _499;
        else
            _500 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _503 <= _502;
        else
            _503 <= _500;
    end
    always @(posedge _84) begin
        if (_82)
            _506 <= _505;
        else
            _506 <= _503;
    end
    always @(posedge _84) begin
        if (_82)
            _509 <= _508;
        else
            _509 <= _506;
    end
    always @(posedge _84) begin
        if (_82)
            _512 <= _511;
        else
            _512 <= _509;
    end
    always @(posedge _84) begin
        if (_82)
            _515 <= _514;
        else
            _515 <= _512;
    end
    always @(posedge _84) begin
        if (_82)
            _518 <= _517;
        else
            _518 <= _515;
    end
    always @(posedge _84) begin
        if (_82)
            _521 <= _520;
        else
            _521 <= _518;
    end
    always @(posedge _84) begin
        if (_82)
            _524 <= _523;
        else
            _524 <= _521;
    end
    assign _553 = _524 & _552;
    assign _554 = _129 & _553;
    assign write_enable_22 = _554 & PHASE_4;
    assign _559 = write_enable_22 | read_enable_18;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_10
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_559), .regcea(vdd), .wea(write_enable_22), .addra(address_22), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_13), .regceb(vdd), .web(write_enable_13), .addrb(address_13), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_566[131:131]), .sbiterrb(_566[130:130]), .doutb(_566[129:66]), .dbiterra(_566[65:65]), .sbiterra(_566[64:64]), .douta(_566[63:0]) );
    assign _567 = _566[63:0];
    assign _497 = ~ PHASE_4;
    assign _15 = _497;
    always @(posedge _84) begin
        if (_82)
            PHASE_4 <= _495;
        else
            if (_72)
                PHASE_4 <= _15;
    end
    assign _579 = PHASE_4 ? _578 : _567;
    assign address_23 = _764 ? _199 : _759;
    assign write_enable_23 = _757 & _764;
    assign address_24 = _764 ? _164 : _68;
    assign _766 = ~ _764;
    assign read_enable_19 = _752 & _766;
    assign _764 = ~ PHASE_7;
    assign write_enable_24 = _750 & _764;
    assign _768 = write_enable_24 | read_enable_19;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_11
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_768), .regcea(vdd), .wea(write_enable_24), .addra(address_24), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_23), .regceb(vdd), .web(write_enable_23), .addrb(address_23), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_773[131:131]), .sbiterrb(_773[130:130]), .doutb(_773[129:66]), .dbiterra(_773[65:65]), .sbiterra(_773[64:64]), .douta(_773[63:0]) );
    assign _774 = _773[63:0];
    assign address_25 = PHASE_7 ? _199 : _759;
    assign _757 = _129 & _720;
    assign write_enable_25 = _757 & PHASE_7;
    assign _682 = _674[129:66];
    assign _681 = _661[129:66];
    assign _683 = PHASE_5 ? _682 : _681;
    assign _679 = _619[129:66];
    assign _678 = _605[129:66];
    assign q1_1 = PHASE_6 ? _679 : _678;
    assign _684 = _586 ? _683 : q1_1;
    assign address_26 = _663 ? _657 : _656;
    assign _669 = ~ _663;
    assign read_enable_20 = _102 & _669;
    assign address_27 = _663 ? _60 : _639;
    assign _665 = ~ _663;
    assign read_enable_21 = _102 & _665;
    assign _663 = ~ PHASE_5;
    assign write_enable_27 = _622 & _663;
    assign _667 = write_enable_27 | read_enable_21;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_12
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_667), .regcea(vdd), .wea(write_enable_27), .addra(address_27), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_20), .regceb(vdd), .web(write_enable_26), .addrb(address_26), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_674[131:131]), .sbiterrb(_674[130:130]), .doutb(_674[129:66]), .dbiterra(_674[65:65]), .sbiterra(_674[64:64]), .douta(_674[63:0]) );
    assign _675 = _674[63:0];
    assign _655 = _172[11:11];
    assign _654 = _172[10:10];
    assign _653 = _172[9:9];
    assign _652 = _172[8:8];
    assign _651 = _172[7:7];
    assign _650 = _172[6:6];
    assign _649 = _172[5:5];
    assign _648 = _172[4:4];
    assign _647 = _172[3:3];
    assign _646 = _172[2:2];
    assign _645 = _172[1:1];
    assign _644 = _172[0:0];
    assign _656 = { _644, _645, _646, _647, _648, _649, _650, _651, _652, _653, _654, _655 };
    assign address_28 = PHASE_5 ? _657 : _656;
    assign _641 = ~ PHASE_5;
    assign read_enable_22 = _102 & _641;
    assign data_25 = wr_d5;
    assign _638 = _137[11:11];
    assign _637 = _137[10:10];
    assign _636 = _137[9:9];
    assign _635 = _137[8:8];
    assign _634 = _137[7:7];
    assign _633 = _137[6:6];
    assign _632 = _137[5:5];
    assign _631 = _137[4:4];
    assign _630 = _137[3:3];
    assign _629 = _137[2:2];
    assign _628 = _137[1:1];
    assign _627 = _137[0:0];
    assign _639 = { _627, _628, _629, _630, _631, _632, _633, _634, _635, _636, _637, _638 };
    assign address_29 = PHASE_5 ? _60 : _639;
    assign _624 = ~ PHASE_5;
    assign read_enable_23 = _102 & _624;
    assign _622 = _62[5:5];
    assign write_enable_29 = _622 & PHASE_5;
    assign _626 = write_enable_29 | read_enable_23;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_13
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_626), .regcea(vdd), .wea(write_enable_29), .addra(address_29), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_22), .regceb(vdd), .web(write_enable_28), .addrb(address_28), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_661[131:131]), .sbiterrb(_661[130:130]), .doutb(_661[129:66]), .dbiterra(_661[65:65]), .sbiterra(_661[64:64]), .douta(_661[63:0]) );
    assign _662 = _661[63:0];
    assign _583 = ~ PHASE_5;
    assign _19 = _583;
    always @(posedge _84) begin
        if (_82)
            PHASE_5 <= _581;
        else
            if (_72)
                PHASE_5 <= _19;
    end
    assign _676 = PHASE_5 ? _675 : _662;
    assign address_30 = _607 ? _199 : _172;
    assign _614 = ~ _607;
    assign read_enable_24 = _102 & _614;
    assign write_enable_30 = _598 & _607;
    assign _616 = write_enable_30 | read_enable_24;
    assign address_31 = _607 ? _164 : _137;
    assign _609 = ~ _607;
    assign read_enable_25 = _102 & _609;
    assign _607 = ~ PHASE_6;
    assign write_enable_31 = _591 & _607;
    assign _611 = write_enable_31 | read_enable_25;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_14
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_611), .regcea(vdd), .wea(write_enable_31), .addra(address_31), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_616), .regceb(vdd), .web(write_enable_30), .addrb(address_30), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_619[131:131]), .sbiterrb(_619[130:130]), .doutb(_619[129:66]), .dbiterra(_619[65:65]), .sbiterra(_619[64:64]), .douta(_619[63:0]) );
    assign _620 = _619[63:0];
    assign _687 = _686[127:64];
    assign data_27 = _687;
    assign address_32 = PHASE_6 ? _199 : _172;
    assign _600 = ~ PHASE_6;
    assign read_enable_26 = _102 & _600;
    assign _597 = ~ _130;
    assign _598 = _129 & _597;
    assign write_enable_32 = _598 & PHASE_6;
    assign _602 = write_enable_32 | read_enable_26;
    assign address_33 = PHASE_6 ? _164 : _137;
    assign _593 = ~ PHASE_6;
    assign read_enable_27 = _102 & _593;
    assign _590 = ~ _130;
    assign _591 = _129 & _590;
    assign write_enable_33 = _591 & PHASE_6;
    assign _595 = write_enable_33 | read_enable_27;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_15
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_595), .regcea(vdd), .wea(write_enable_33), .addra(address_33), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_602), .regceb(vdd), .web(write_enable_32), .addrb(address_32), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_605[131:131]), .sbiterrb(_605[130:130]), .doutb(_605[129:66]), .dbiterra(_605[65:65]), .sbiterra(_605[64:64]), .douta(_605[63:0]) );
    assign _606 = _605[63:0];
    assign _688 = ~ PHASE_6;
    assign _21 = _688;
    always @(posedge _84) begin
        if (_82)
            PHASE_6 <= _588;
        else
            if (_99)
                PHASE_6 <= _21;
    end
    assign q0_1 = PHASE_6 ? _620 : _606;
    always @(posedge _84) begin
        if (_82)
            _586 <= _585;
        else
            _586 <= _92;
    end
    assign _677 = _586 ? _676 : q0_1;
    dp_52
        dp_4
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_677), .d2(_684), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_686[191:128]), .q2(_686[127:64]), .q1(_686[63:0]) );
    assign _689 = _686[63:0];
    assign data_31 = _689;
    assign address_34 = PHASE_7 ? _164 : _68;
    assign _753 = ~ PHASE_7;
    assign _752 = _70[5:5];
    assign read_enable_28 = _752 & _753;
    always @(posedge _84) begin
        if (_82)
            _723 <= _722;
        else
            _723 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _726 <= _725;
        else
            _726 <= _723;
    end
    always @(posedge _84) begin
        if (_82)
            _729 <= _728;
        else
            _729 <= _726;
    end
    always @(posedge _84) begin
        if (_82)
            _732 <= _731;
        else
            _732 <= _729;
    end
    always @(posedge _84) begin
        if (_82)
            _735 <= _734;
        else
            _735 <= _732;
    end
    always @(posedge _84) begin
        if (_82)
            _738 <= _737;
        else
            _738 <= _735;
    end
    always @(posedge _84) begin
        if (_82)
            _741 <= _740;
        else
            _741 <= _738;
    end
    always @(posedge _84) begin
        if (_82)
            _744 <= _743;
        else
            _744 <= _741;
    end
    always @(posedge _84) begin
        if (_82)
            _747 <= _746;
        else
            _747 <= _744;
    end
    assign _748 = ~ _747;
    always @(posedge _84) begin
        if (_82)
            _696 <= _695;
        else
            _696 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _699 <= _698;
        else
            _699 <= _696;
    end
    always @(posedge _84) begin
        if (_82)
            _702 <= _701;
        else
            _702 <= _699;
    end
    always @(posedge _84) begin
        if (_82)
            _705 <= _704;
        else
            _705 <= _702;
    end
    always @(posedge _84) begin
        if (_82)
            _708 <= _707;
        else
            _708 <= _705;
    end
    always @(posedge _84) begin
        if (_82)
            _711 <= _710;
        else
            _711 <= _708;
    end
    always @(posedge _84) begin
        if (_82)
            _714 <= _713;
        else
            _714 <= _711;
    end
    always @(posedge _84) begin
        if (_82)
            _717 <= _716;
        else
            _717 <= _714;
    end
    always @(posedge _84) begin
        if (_82)
            _720 <= _719;
        else
            _720 <= _717;
    end
    assign _749 = _720 & _748;
    assign _750 = _129 & _749;
    assign write_enable_34 = _750 & PHASE_7;
    assign _755 = write_enable_34 | read_enable_28;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_16
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_755), .regcea(vdd), .wea(write_enable_34), .addra(address_34), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_25), .regceb(vdd), .web(write_enable_25), .addrb(address_25), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_762[131:131]), .sbiterrb(_762[130:130]), .doutb(_762[129:66]), .dbiterra(_762[65:65]), .sbiterra(_762[64:64]), .douta(_762[63:0]) );
    assign _763 = _762[63:0];
    assign _693 = ~ PHASE_7;
    assign _23 = _693;
    always @(posedge _84) begin
        if (_82)
            PHASE_7 <= _691;
        else
            if (_72)
                PHASE_7 <= _23;
    end
    assign _775 = PHASE_7 ? _774 : _763;
    assign address_35 = _960 ? _199 : _955;
    assign write_enable_35 = _953 & _960;
    assign address_36 = _960 ? _164 : _68;
    assign _962 = ~ _960;
    assign read_enable_29 = _948 & _962;
    assign _960 = ~ PHASE_10;
    assign write_enable_36 = _946 & _960;
    assign _964 = write_enable_36 | read_enable_29;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_17
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_964), .regcea(vdd), .wea(write_enable_36), .addra(address_36), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_35), .regceb(vdd), .web(write_enable_35), .addrb(address_35), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_969[131:131]), .sbiterrb(_969[130:130]), .doutb(_969[129:66]), .dbiterra(_969[65:65]), .sbiterra(_969[64:64]), .douta(_969[63:0]) );
    assign _970 = _969[63:0];
    assign address_37 = PHASE_10 ? _199 : _955;
    assign _953 = _129 & _916;
    assign write_enable_37 = _953 & PHASE_10;
    assign _878 = _870[129:66];
    assign _877 = _857[129:66];
    assign _879 = PHASE_8 ? _878 : _877;
    assign _875 = _815[129:66];
    assign _874 = _801[129:66];
    assign q1_2 = PHASE_9 ? _875 : _874;
    assign _880 = _782 ? _879 : q1_2;
    assign address_38 = _859 ? _853 : _852;
    assign _865 = ~ _859;
    assign read_enable_30 = _102 & _865;
    assign address_39 = _859 ? _60 : _835;
    assign _861 = ~ _859;
    assign read_enable_31 = _102 & _861;
    assign _859 = ~ PHASE_8;
    assign write_enable_39 = _818 & _859;
    assign _863 = write_enable_39 | read_enable_31;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_18
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_863), .regcea(vdd), .wea(write_enable_39), .addra(address_39), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_30), .regceb(vdd), .web(write_enable_38), .addrb(address_38), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_870[131:131]), .sbiterrb(_870[130:130]), .doutb(_870[129:66]), .dbiterra(_870[65:65]), .sbiterra(_870[64:64]), .douta(_870[63:0]) );
    assign _871 = _870[63:0];
    assign _851 = _172[11:11];
    assign _850 = _172[10:10];
    assign _849 = _172[9:9];
    assign _848 = _172[8:8];
    assign _847 = _172[7:7];
    assign _846 = _172[6:6];
    assign _845 = _172[5:5];
    assign _844 = _172[4:4];
    assign _843 = _172[3:3];
    assign _842 = _172[2:2];
    assign _841 = _172[1:1];
    assign _840 = _172[0:0];
    assign _852 = { _840, _841, _842, _843, _844, _845, _846, _847, _848, _849, _850, _851 };
    assign address_40 = PHASE_8 ? _853 : _852;
    assign _837 = ~ PHASE_8;
    assign read_enable_32 = _102 & _837;
    assign data_37 = wr_d4;
    assign _834 = _137[11:11];
    assign _833 = _137[10:10];
    assign _832 = _137[9:9];
    assign _831 = _137[8:8];
    assign _830 = _137[7:7];
    assign _829 = _137[6:6];
    assign _828 = _137[5:5];
    assign _827 = _137[4:4];
    assign _826 = _137[3:3];
    assign _825 = _137[2:2];
    assign _824 = _137[1:1];
    assign _823 = _137[0:0];
    assign _835 = { _823, _824, _825, _826, _827, _828, _829, _830, _831, _832, _833, _834 };
    assign address_41 = PHASE_8 ? _60 : _835;
    assign _820 = ~ PHASE_8;
    assign read_enable_33 = _102 & _820;
    assign _818 = _62[4:4];
    assign write_enable_41 = _818 & PHASE_8;
    assign _822 = write_enable_41 | read_enable_33;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_19
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_822), .regcea(vdd), .wea(write_enable_41), .addra(address_41), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_32), .regceb(vdd), .web(write_enable_40), .addrb(address_40), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_857[131:131]), .sbiterrb(_857[130:130]), .doutb(_857[129:66]), .dbiterra(_857[65:65]), .sbiterra(_857[64:64]), .douta(_857[63:0]) );
    assign _858 = _857[63:0];
    assign _779 = ~ PHASE_8;
    assign _27 = _779;
    always @(posedge _84) begin
        if (_82)
            PHASE_8 <= _777;
        else
            if (_72)
                PHASE_8 <= _27;
    end
    assign _872 = PHASE_8 ? _871 : _858;
    assign address_42 = _803 ? _199 : _172;
    assign _810 = ~ _803;
    assign read_enable_34 = _102 & _810;
    assign write_enable_42 = _794 & _803;
    assign _812 = write_enable_42 | read_enable_34;
    assign address_43 = _803 ? _164 : _137;
    assign _805 = ~ _803;
    assign read_enable_35 = _102 & _805;
    assign _803 = ~ PHASE_9;
    assign write_enable_43 = _787 & _803;
    assign _807 = write_enable_43 | read_enable_35;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_20
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_807), .regcea(vdd), .wea(write_enable_43), .addra(address_43), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_812), .regceb(vdd), .web(write_enable_42), .addrb(address_42), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_815[131:131]), .sbiterrb(_815[130:130]), .doutb(_815[129:66]), .dbiterra(_815[65:65]), .sbiterra(_815[64:64]), .douta(_815[63:0]) );
    assign _816 = _815[63:0];
    assign _883 = _882[127:64];
    assign data_39 = _883;
    assign address_44 = PHASE_9 ? _199 : _172;
    assign _796 = ~ PHASE_9;
    assign read_enable_36 = _102 & _796;
    assign _793 = ~ _130;
    assign _794 = _129 & _793;
    assign write_enable_44 = _794 & PHASE_9;
    assign _798 = write_enable_44 | read_enable_36;
    assign address_45 = PHASE_9 ? _164 : _137;
    assign _789 = ~ PHASE_9;
    assign read_enable_37 = _102 & _789;
    assign _786 = ~ _130;
    assign _787 = _129 & _786;
    assign write_enable_45 = _787 & PHASE_9;
    assign _791 = write_enable_45 | read_enable_37;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_21
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_791), .regcea(vdd), .wea(write_enable_45), .addra(address_45), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_798), .regceb(vdd), .web(write_enable_44), .addrb(address_44), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_801[131:131]), .sbiterrb(_801[130:130]), .doutb(_801[129:66]), .dbiterra(_801[65:65]), .sbiterra(_801[64:64]), .douta(_801[63:0]) );
    assign _802 = _801[63:0];
    assign _884 = ~ PHASE_9;
    assign _29 = _884;
    always @(posedge _84) begin
        if (_82)
            PHASE_9 <= _784;
        else
            if (_99)
                PHASE_9 <= _29;
    end
    assign q0_2 = PHASE_9 ? _816 : _802;
    always @(posedge _84) begin
        if (_82)
            _782 <= _781;
        else
            _782 <= _92;
    end
    assign _873 = _782 ? _872 : q0_2;
    dp_51
        dp_3
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_873), .d2(_880), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_882[191:128]), .q2(_882[127:64]), .q1(_882[63:0]) );
    assign _885 = _882[63:0];
    assign data_43 = _885;
    assign address_46 = PHASE_10 ? _164 : _68;
    assign _949 = ~ PHASE_10;
    assign _948 = _70[4:4];
    assign read_enable_38 = _948 & _949;
    always @(posedge _84) begin
        if (_82)
            _919 <= _918;
        else
            _919 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _922 <= _921;
        else
            _922 <= _919;
    end
    always @(posedge _84) begin
        if (_82)
            _925 <= _924;
        else
            _925 <= _922;
    end
    always @(posedge _84) begin
        if (_82)
            _928 <= _927;
        else
            _928 <= _925;
    end
    always @(posedge _84) begin
        if (_82)
            _931 <= _930;
        else
            _931 <= _928;
    end
    always @(posedge _84) begin
        if (_82)
            _934 <= _933;
        else
            _934 <= _931;
    end
    always @(posedge _84) begin
        if (_82)
            _937 <= _936;
        else
            _937 <= _934;
    end
    always @(posedge _84) begin
        if (_82)
            _940 <= _939;
        else
            _940 <= _937;
    end
    always @(posedge _84) begin
        if (_82)
            _943 <= _942;
        else
            _943 <= _940;
    end
    assign _944 = ~ _943;
    always @(posedge _84) begin
        if (_82)
            _892 <= _891;
        else
            _892 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _895 <= _894;
        else
            _895 <= _892;
    end
    always @(posedge _84) begin
        if (_82)
            _898 <= _897;
        else
            _898 <= _895;
    end
    always @(posedge _84) begin
        if (_82)
            _901 <= _900;
        else
            _901 <= _898;
    end
    always @(posedge _84) begin
        if (_82)
            _904 <= _903;
        else
            _904 <= _901;
    end
    always @(posedge _84) begin
        if (_82)
            _907 <= _906;
        else
            _907 <= _904;
    end
    always @(posedge _84) begin
        if (_82)
            _910 <= _909;
        else
            _910 <= _907;
    end
    always @(posedge _84) begin
        if (_82)
            _913 <= _912;
        else
            _913 <= _910;
    end
    always @(posedge _84) begin
        if (_82)
            _916 <= _915;
        else
            _916 <= _913;
    end
    assign _945 = _916 & _944;
    assign _946 = _129 & _945;
    assign write_enable_46 = _946 & PHASE_10;
    assign _951 = write_enable_46 | read_enable_38;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_22
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_951), .regcea(vdd), .wea(write_enable_46), .addra(address_46), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_37), .regceb(vdd), .web(write_enable_37), .addrb(address_37), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_958[131:131]), .sbiterrb(_958[130:130]), .doutb(_958[129:66]), .dbiterra(_958[65:65]), .sbiterra(_958[64:64]), .douta(_958[63:0]) );
    assign _959 = _958[63:0];
    assign _889 = ~ PHASE_10;
    assign _31 = _889;
    always @(posedge _84) begin
        if (_82)
            PHASE_10 <= _887;
        else
            if (_72)
                PHASE_10 <= _31;
    end
    assign _971 = PHASE_10 ? _970 : _959;
    assign address_47 = _1156 ? _199 : _1151;
    assign write_enable_47 = _1149 & _1156;
    assign address_48 = _1156 ? _164 : _68;
    assign _1158 = ~ _1156;
    assign read_enable_39 = _1144 & _1158;
    assign _1156 = ~ PHASE_13;
    assign write_enable_48 = _1142 & _1156;
    assign _1160 = write_enable_48 | read_enable_39;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_23
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1160), .regcea(vdd), .wea(write_enable_48), .addra(address_48), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_47), .regceb(vdd), .web(write_enable_47), .addrb(address_47), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1165[131:131]), .sbiterrb(_1165[130:130]), .doutb(_1165[129:66]), .dbiterra(_1165[65:65]), .sbiterra(_1165[64:64]), .douta(_1165[63:0]) );
    assign _1166 = _1165[63:0];
    assign address_49 = PHASE_13 ? _199 : _1151;
    assign _1149 = _129 & _1112;
    assign write_enable_49 = _1149 & PHASE_13;
    assign _1074 = _1066[129:66];
    assign _1073 = _1053[129:66];
    assign _1075 = PHASE_11 ? _1074 : _1073;
    assign _1071 = _1011[129:66];
    assign _1070 = _997[129:66];
    assign q1_3 = PHASE_12 ? _1071 : _1070;
    assign _1076 = _978 ? _1075 : q1_3;
    assign address_50 = _1055 ? _1049 : _1048;
    assign _1061 = ~ _1055;
    assign read_enable_40 = _102 & _1061;
    assign address_51 = _1055 ? _60 : _1031;
    assign _1057 = ~ _1055;
    assign read_enable_41 = _102 & _1057;
    assign _1055 = ~ PHASE_11;
    assign write_enable_51 = _1014 & _1055;
    assign _1059 = write_enable_51 | read_enable_41;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_24
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1059), .regcea(vdd), .wea(write_enable_51), .addra(address_51), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_40), .regceb(vdd), .web(write_enable_50), .addrb(address_50), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1066[131:131]), .sbiterrb(_1066[130:130]), .doutb(_1066[129:66]), .dbiterra(_1066[65:65]), .sbiterra(_1066[64:64]), .douta(_1066[63:0]) );
    assign _1067 = _1066[63:0];
    assign _1047 = _172[11:11];
    assign _1046 = _172[10:10];
    assign _1045 = _172[9:9];
    assign _1044 = _172[8:8];
    assign _1043 = _172[7:7];
    assign _1042 = _172[6:6];
    assign _1041 = _172[5:5];
    assign _1040 = _172[4:4];
    assign _1039 = _172[3:3];
    assign _1038 = _172[2:2];
    assign _1037 = _172[1:1];
    assign _1036 = _172[0:0];
    assign _1048 = { _1036, _1037, _1038, _1039, _1040, _1041, _1042, _1043, _1044, _1045, _1046, _1047 };
    assign address_52 = PHASE_11 ? _1049 : _1048;
    assign _1033 = ~ PHASE_11;
    assign read_enable_42 = _102 & _1033;
    assign data_49 = wr_d3;
    assign _1030 = _137[11:11];
    assign _1029 = _137[10:10];
    assign _1028 = _137[9:9];
    assign _1027 = _137[8:8];
    assign _1026 = _137[7:7];
    assign _1025 = _137[6:6];
    assign _1024 = _137[5:5];
    assign _1023 = _137[4:4];
    assign _1022 = _137[3:3];
    assign _1021 = _137[2:2];
    assign _1020 = _137[1:1];
    assign _1019 = _137[0:0];
    assign _1031 = { _1019, _1020, _1021, _1022, _1023, _1024, _1025, _1026, _1027, _1028, _1029, _1030 };
    assign address_53 = PHASE_11 ? _60 : _1031;
    assign _1016 = ~ PHASE_11;
    assign read_enable_43 = _102 & _1016;
    assign _1014 = _62[3:3];
    assign write_enable_53 = _1014 & PHASE_11;
    assign _1018 = write_enable_53 | read_enable_43;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_25
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1018), .regcea(vdd), .wea(write_enable_53), .addra(address_53), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_42), .regceb(vdd), .web(write_enable_52), .addrb(address_52), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1053[131:131]), .sbiterrb(_1053[130:130]), .doutb(_1053[129:66]), .dbiterra(_1053[65:65]), .sbiterra(_1053[64:64]), .douta(_1053[63:0]) );
    assign _1054 = _1053[63:0];
    assign _975 = ~ PHASE_11;
    assign _35 = _975;
    always @(posedge _84) begin
        if (_82)
            PHASE_11 <= _973;
        else
            if (_72)
                PHASE_11 <= _35;
    end
    assign _1068 = PHASE_11 ? _1067 : _1054;
    assign address_54 = _999 ? _199 : _172;
    assign _1006 = ~ _999;
    assign read_enable_44 = _102 & _1006;
    assign write_enable_54 = _990 & _999;
    assign _1008 = write_enable_54 | read_enable_44;
    assign address_55 = _999 ? _164 : _137;
    assign _1001 = ~ _999;
    assign read_enable_45 = _102 & _1001;
    assign _999 = ~ PHASE_12;
    assign write_enable_55 = _983 & _999;
    assign _1003 = write_enable_55 | read_enable_45;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_26
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1003), .regcea(vdd), .wea(write_enable_55), .addra(address_55), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1008), .regceb(vdd), .web(write_enable_54), .addrb(address_54), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1011[131:131]), .sbiterrb(_1011[130:130]), .doutb(_1011[129:66]), .dbiterra(_1011[65:65]), .sbiterra(_1011[64:64]), .douta(_1011[63:0]) );
    assign _1012 = _1011[63:0];
    assign _1079 = _1078[127:64];
    assign data_51 = _1079;
    assign address_56 = PHASE_12 ? _199 : _172;
    assign _992 = ~ PHASE_12;
    assign read_enable_46 = _102 & _992;
    assign _989 = ~ _130;
    assign _990 = _129 & _989;
    assign write_enable_56 = _990 & PHASE_12;
    assign _994 = write_enable_56 | read_enable_46;
    assign address_57 = PHASE_12 ? _164 : _137;
    assign _985 = ~ PHASE_12;
    assign read_enable_47 = _102 & _985;
    assign _982 = ~ _130;
    assign _983 = _129 & _982;
    assign write_enable_57 = _983 & PHASE_12;
    assign _987 = write_enable_57 | read_enable_47;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_27
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_987), .regcea(vdd), .wea(write_enable_57), .addra(address_57), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_994), .regceb(vdd), .web(write_enable_56), .addrb(address_56), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_997[131:131]), .sbiterrb(_997[130:130]), .doutb(_997[129:66]), .dbiterra(_997[65:65]), .sbiterra(_997[64:64]), .douta(_997[63:0]) );
    assign _998 = _997[63:0];
    assign _1080 = ~ PHASE_12;
    assign _37 = _1080;
    always @(posedge _84) begin
        if (_82)
            PHASE_12 <= _980;
        else
            if (_99)
                PHASE_12 <= _37;
    end
    assign q0_3 = PHASE_12 ? _1012 : _998;
    always @(posedge _84) begin
        if (_82)
            _978 <= _977;
        else
            _978 <= _92;
    end
    assign _1069 = _978 ? _1068 : q0_3;
    dp_50
        dp_2
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1069), .d2(_1076), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1078[191:128]), .q2(_1078[127:64]), .q1(_1078[63:0]) );
    assign _1081 = _1078[63:0];
    assign data_55 = _1081;
    assign address_58 = PHASE_13 ? _164 : _68;
    assign _1145 = ~ PHASE_13;
    assign _1144 = _70[3:3];
    assign read_enable_48 = _1144 & _1145;
    always @(posedge _84) begin
        if (_82)
            _1115 <= _1114;
        else
            _1115 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1118 <= _1117;
        else
            _1118 <= _1115;
    end
    always @(posedge _84) begin
        if (_82)
            _1121 <= _1120;
        else
            _1121 <= _1118;
    end
    always @(posedge _84) begin
        if (_82)
            _1124 <= _1123;
        else
            _1124 <= _1121;
    end
    always @(posedge _84) begin
        if (_82)
            _1127 <= _1126;
        else
            _1127 <= _1124;
    end
    always @(posedge _84) begin
        if (_82)
            _1130 <= _1129;
        else
            _1130 <= _1127;
    end
    always @(posedge _84) begin
        if (_82)
            _1133 <= _1132;
        else
            _1133 <= _1130;
    end
    always @(posedge _84) begin
        if (_82)
            _1136 <= _1135;
        else
            _1136 <= _1133;
    end
    always @(posedge _84) begin
        if (_82)
            _1139 <= _1138;
        else
            _1139 <= _1136;
    end
    assign _1140 = ~ _1139;
    always @(posedge _84) begin
        if (_82)
            _1088 <= _1087;
        else
            _1088 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1091 <= _1090;
        else
            _1091 <= _1088;
    end
    always @(posedge _84) begin
        if (_82)
            _1094 <= _1093;
        else
            _1094 <= _1091;
    end
    always @(posedge _84) begin
        if (_82)
            _1097 <= _1096;
        else
            _1097 <= _1094;
    end
    always @(posedge _84) begin
        if (_82)
            _1100 <= _1099;
        else
            _1100 <= _1097;
    end
    always @(posedge _84) begin
        if (_82)
            _1103 <= _1102;
        else
            _1103 <= _1100;
    end
    always @(posedge _84) begin
        if (_82)
            _1106 <= _1105;
        else
            _1106 <= _1103;
    end
    always @(posedge _84) begin
        if (_82)
            _1109 <= _1108;
        else
            _1109 <= _1106;
    end
    always @(posedge _84) begin
        if (_82)
            _1112 <= _1111;
        else
            _1112 <= _1109;
    end
    assign _1141 = _1112 & _1140;
    assign _1142 = _129 & _1141;
    assign write_enable_58 = _1142 & PHASE_13;
    assign _1147 = write_enable_58 | read_enable_48;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_28
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1147), .regcea(vdd), .wea(write_enable_58), .addra(address_58), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_49), .regceb(vdd), .web(write_enable_49), .addrb(address_49), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1154[131:131]), .sbiterrb(_1154[130:130]), .doutb(_1154[129:66]), .dbiterra(_1154[65:65]), .sbiterra(_1154[64:64]), .douta(_1154[63:0]) );
    assign _1155 = _1154[63:0];
    assign _1085 = ~ PHASE_13;
    assign _39 = _1085;
    always @(posedge _84) begin
        if (_82)
            PHASE_13 <= _1083;
        else
            if (_72)
                PHASE_13 <= _39;
    end
    assign _1167 = PHASE_13 ? _1166 : _1155;
    assign address_59 = _1352 ? _199 : _1347;
    assign write_enable_59 = _1345 & _1352;
    assign address_60 = _1352 ? _164 : _68;
    assign _1354 = ~ _1352;
    assign read_enable_49 = _1340 & _1354;
    assign _1352 = ~ PHASE_16;
    assign write_enable_60 = _1338 & _1352;
    assign _1356 = write_enable_60 | read_enable_49;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_29
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1356), .regcea(vdd), .wea(write_enable_60), .addra(address_60), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_59), .regceb(vdd), .web(write_enable_59), .addrb(address_59), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1361[131:131]), .sbiterrb(_1361[130:130]), .doutb(_1361[129:66]), .dbiterra(_1361[65:65]), .sbiterra(_1361[64:64]), .douta(_1361[63:0]) );
    assign _1362 = _1361[63:0];
    assign address_61 = PHASE_16 ? _199 : _1347;
    assign _1345 = _129 & _1308;
    assign write_enable_61 = _1345 & PHASE_16;
    assign _1270 = _1262[129:66];
    assign _1269 = _1249[129:66];
    assign _1271 = PHASE_14 ? _1270 : _1269;
    assign _1267 = _1207[129:66];
    assign _1266 = _1193[129:66];
    assign q1_4 = PHASE_15 ? _1267 : _1266;
    assign _1272 = _1174 ? _1271 : q1_4;
    assign address_62 = _1251 ? _1245 : _1244;
    assign _1257 = ~ _1251;
    assign read_enable_50 = _102 & _1257;
    assign address_63 = _1251 ? _60 : _1227;
    assign _1253 = ~ _1251;
    assign read_enable_51 = _102 & _1253;
    assign _1251 = ~ PHASE_14;
    assign write_enable_63 = _1210 & _1251;
    assign _1255 = write_enable_63 | read_enable_51;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_30
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1255), .regcea(vdd), .wea(write_enable_63), .addra(address_63), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_50), .regceb(vdd), .web(write_enable_62), .addrb(address_62), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1262[131:131]), .sbiterrb(_1262[130:130]), .doutb(_1262[129:66]), .dbiterra(_1262[65:65]), .sbiterra(_1262[64:64]), .douta(_1262[63:0]) );
    assign _1263 = _1262[63:0];
    assign _1243 = _172[11:11];
    assign _1242 = _172[10:10];
    assign _1241 = _172[9:9];
    assign _1240 = _172[8:8];
    assign _1239 = _172[7:7];
    assign _1238 = _172[6:6];
    assign _1237 = _172[5:5];
    assign _1236 = _172[4:4];
    assign _1235 = _172[3:3];
    assign _1234 = _172[2:2];
    assign _1233 = _172[1:1];
    assign _1232 = _172[0:0];
    assign _1244 = { _1232, _1233, _1234, _1235, _1236, _1237, _1238, _1239, _1240, _1241, _1242, _1243 };
    assign address_64 = PHASE_14 ? _1245 : _1244;
    assign _1229 = ~ PHASE_14;
    assign read_enable_52 = _102 & _1229;
    assign data_61 = wr_d2;
    assign _1226 = _137[11:11];
    assign _1225 = _137[10:10];
    assign _1224 = _137[9:9];
    assign _1223 = _137[8:8];
    assign _1222 = _137[7:7];
    assign _1221 = _137[6:6];
    assign _1220 = _137[5:5];
    assign _1219 = _137[4:4];
    assign _1218 = _137[3:3];
    assign _1217 = _137[2:2];
    assign _1216 = _137[1:1];
    assign _1215 = _137[0:0];
    assign _1227 = { _1215, _1216, _1217, _1218, _1219, _1220, _1221, _1222, _1223, _1224, _1225, _1226 };
    assign address_65 = PHASE_14 ? _60 : _1227;
    assign _1212 = ~ PHASE_14;
    assign read_enable_53 = _102 & _1212;
    assign _1210 = _62[2:2];
    assign write_enable_65 = _1210 & PHASE_14;
    assign _1214 = write_enable_65 | read_enable_53;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_31
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1214), .regcea(vdd), .wea(write_enable_65), .addra(address_65), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_52), .regceb(vdd), .web(write_enable_64), .addrb(address_64), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1249[131:131]), .sbiterrb(_1249[130:130]), .doutb(_1249[129:66]), .dbiterra(_1249[65:65]), .sbiterra(_1249[64:64]), .douta(_1249[63:0]) );
    assign _1250 = _1249[63:0];
    assign _1171 = ~ PHASE_14;
    assign _43 = _1171;
    always @(posedge _84) begin
        if (_82)
            PHASE_14 <= _1169;
        else
            if (_72)
                PHASE_14 <= _43;
    end
    assign _1264 = PHASE_14 ? _1263 : _1250;
    assign address_66 = _1195 ? _199 : _172;
    assign _1202 = ~ _1195;
    assign read_enable_54 = _102 & _1202;
    assign write_enable_66 = _1186 & _1195;
    assign _1204 = write_enable_66 | read_enable_54;
    assign address_67 = _1195 ? _164 : _137;
    assign _1197 = ~ _1195;
    assign read_enable_55 = _102 & _1197;
    assign _1195 = ~ PHASE_15;
    assign write_enable_67 = _1179 & _1195;
    assign _1199 = write_enable_67 | read_enable_55;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_32
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1199), .regcea(vdd), .wea(write_enable_67), .addra(address_67), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1204), .regceb(vdd), .web(write_enable_66), .addrb(address_66), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1207[131:131]), .sbiterrb(_1207[130:130]), .doutb(_1207[129:66]), .dbiterra(_1207[65:65]), .sbiterra(_1207[64:64]), .douta(_1207[63:0]) );
    assign _1208 = _1207[63:0];
    assign _1275 = _1274[127:64];
    assign data_63 = _1275;
    assign address_68 = PHASE_15 ? _199 : _172;
    assign _1188 = ~ PHASE_15;
    assign read_enable_56 = _102 & _1188;
    assign _1185 = ~ _130;
    assign _1186 = _129 & _1185;
    assign write_enable_68 = _1186 & PHASE_15;
    assign _1190 = write_enable_68 | read_enable_56;
    assign address_69 = PHASE_15 ? _164 : _137;
    assign _1181 = ~ PHASE_15;
    assign read_enable_57 = _102 & _1181;
    assign _1178 = ~ _130;
    assign _1179 = _129 & _1178;
    assign write_enable_69 = _1179 & PHASE_15;
    assign _1183 = write_enable_69 | read_enable_57;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_33
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1183), .regcea(vdd), .wea(write_enable_69), .addra(address_69), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1190), .regceb(vdd), .web(write_enable_68), .addrb(address_68), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1193[131:131]), .sbiterrb(_1193[130:130]), .doutb(_1193[129:66]), .dbiterra(_1193[65:65]), .sbiterra(_1193[64:64]), .douta(_1193[63:0]) );
    assign _1194 = _1193[63:0];
    assign _1276 = ~ PHASE_15;
    assign _45 = _1276;
    always @(posedge _84) begin
        if (_82)
            PHASE_15 <= _1176;
        else
            if (_99)
                PHASE_15 <= _45;
    end
    assign q0_4 = PHASE_15 ? _1208 : _1194;
    always @(posedge _84) begin
        if (_82)
            _1174 <= _1173;
        else
            _1174 <= _92;
    end
    assign _1265 = _1174 ? _1264 : q0_4;
    dp_49
        dp_1
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1265), .d2(_1272), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1274[191:128]), .q2(_1274[127:64]), .q1(_1274[63:0]) );
    assign _1277 = _1274[63:0];
    assign data_67 = _1277;
    assign address_70 = PHASE_16 ? _164 : _68;
    assign _1341 = ~ PHASE_16;
    assign _1340 = _70[2:2];
    assign read_enable_58 = _1340 & _1341;
    always @(posedge _84) begin
        if (_82)
            _1311 <= _1310;
        else
            _1311 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1314 <= _1313;
        else
            _1314 <= _1311;
    end
    always @(posedge _84) begin
        if (_82)
            _1317 <= _1316;
        else
            _1317 <= _1314;
    end
    always @(posedge _84) begin
        if (_82)
            _1320 <= _1319;
        else
            _1320 <= _1317;
    end
    always @(posedge _84) begin
        if (_82)
            _1323 <= _1322;
        else
            _1323 <= _1320;
    end
    always @(posedge _84) begin
        if (_82)
            _1326 <= _1325;
        else
            _1326 <= _1323;
    end
    always @(posedge _84) begin
        if (_82)
            _1329 <= _1328;
        else
            _1329 <= _1326;
    end
    always @(posedge _84) begin
        if (_82)
            _1332 <= _1331;
        else
            _1332 <= _1329;
    end
    always @(posedge _84) begin
        if (_82)
            _1335 <= _1334;
        else
            _1335 <= _1332;
    end
    assign _1336 = ~ _1335;
    always @(posedge _84) begin
        if (_82)
            _1284 <= _1283;
        else
            _1284 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1287 <= _1286;
        else
            _1287 <= _1284;
    end
    always @(posedge _84) begin
        if (_82)
            _1290 <= _1289;
        else
            _1290 <= _1287;
    end
    always @(posedge _84) begin
        if (_82)
            _1293 <= _1292;
        else
            _1293 <= _1290;
    end
    always @(posedge _84) begin
        if (_82)
            _1296 <= _1295;
        else
            _1296 <= _1293;
    end
    always @(posedge _84) begin
        if (_82)
            _1299 <= _1298;
        else
            _1299 <= _1296;
    end
    always @(posedge _84) begin
        if (_82)
            _1302 <= _1301;
        else
            _1302 <= _1299;
    end
    always @(posedge _84) begin
        if (_82)
            _1305 <= _1304;
        else
            _1305 <= _1302;
    end
    always @(posedge _84) begin
        if (_82)
            _1308 <= _1307;
        else
            _1308 <= _1305;
    end
    assign _1337 = _1308 & _1336;
    assign _1338 = _129 & _1337;
    assign write_enable_70 = _1338 & PHASE_16;
    assign _1343 = write_enable_70 | read_enable_58;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_34
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1343), .regcea(vdd), .wea(write_enable_70), .addra(address_70), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_61), .regceb(vdd), .web(write_enable_61), .addrb(address_61), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1350[131:131]), .sbiterrb(_1350[130:130]), .doutb(_1350[129:66]), .dbiterra(_1350[65:65]), .sbiterra(_1350[64:64]), .douta(_1350[63:0]) );
    assign _1351 = _1350[63:0];
    assign _1281 = ~ PHASE_16;
    assign _47 = _1281;
    always @(posedge _84) begin
        if (_82)
            PHASE_16 <= _1279;
        else
            if (_72)
                PHASE_16 <= _47;
    end
    assign _1363 = PHASE_16 ? _1362 : _1351;
    assign address_71 = _1548 ? _199 : _1543;
    assign write_enable_71 = _1541 & _1548;
    assign address_72 = _1548 ? _164 : _68;
    assign _1550 = ~ _1548;
    assign read_enable_59 = _1536 & _1550;
    assign _1548 = ~ PHASE_19;
    assign write_enable_72 = _1534 & _1548;
    assign _1552 = write_enable_72 | read_enable_59;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_35
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1552), .regcea(vdd), .wea(write_enable_72), .addra(address_72), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_71), .regceb(vdd), .web(write_enable_71), .addrb(address_71), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1557[131:131]), .sbiterrb(_1557[130:130]), .doutb(_1557[129:66]), .dbiterra(_1557[65:65]), .sbiterra(_1557[64:64]), .douta(_1557[63:0]) );
    assign _1558 = _1557[63:0];
    assign address_73 = PHASE_19 ? _199 : _1543;
    assign _1541 = _129 & _1504;
    assign write_enable_73 = _1541 & PHASE_19;
    assign _1466 = _1458[129:66];
    assign _1465 = _1445[129:66];
    assign _1467 = PHASE_17 ? _1466 : _1465;
    assign _1463 = _1403[129:66];
    assign _1462 = _1389[129:66];
    assign q1_5 = PHASE_18 ? _1463 : _1462;
    assign _1468 = _1370 ? _1467 : q1_5;
    assign address_74 = _1447 ? _1441 : _1440;
    assign _1453 = ~ _1447;
    assign read_enable_60 = _102 & _1453;
    assign address_75 = _1447 ? _60 : _1423;
    assign _1449 = ~ _1447;
    assign read_enable_61 = _102 & _1449;
    assign _1447 = ~ PHASE_17;
    assign write_enable_75 = _1406 & _1447;
    assign _1451 = write_enable_75 | read_enable_61;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_36
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1451), .regcea(vdd), .wea(write_enable_75), .addra(address_75), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_60), .regceb(vdd), .web(write_enable_74), .addrb(address_74), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1458[131:131]), .sbiterrb(_1458[130:130]), .doutb(_1458[129:66]), .dbiterra(_1458[65:65]), .sbiterra(_1458[64:64]), .douta(_1458[63:0]) );
    assign _1459 = _1458[63:0];
    assign _1439 = _172[11:11];
    assign _1438 = _172[10:10];
    assign _1437 = _172[9:9];
    assign _1436 = _172[8:8];
    assign _1435 = _172[7:7];
    assign _1434 = _172[6:6];
    assign _1433 = _172[5:5];
    assign _1432 = _172[4:4];
    assign _1431 = _172[3:3];
    assign _1430 = _172[2:2];
    assign _1429 = _172[1:1];
    assign _1428 = _172[0:0];
    assign _1440 = { _1428, _1429, _1430, _1431, _1432, _1433, _1434, _1435, _1436, _1437, _1438, _1439 };
    assign address_76 = PHASE_17 ? _1441 : _1440;
    assign _1425 = ~ PHASE_17;
    assign read_enable_62 = _102 & _1425;
    assign data_73 = wr_d1;
    assign _1422 = _137[11:11];
    assign _1421 = _137[10:10];
    assign _1420 = _137[9:9];
    assign _1419 = _137[8:8];
    assign _1418 = _137[7:7];
    assign _1417 = _137[6:6];
    assign _1416 = _137[5:5];
    assign _1415 = _137[4:4];
    assign _1414 = _137[3:3];
    assign _1413 = _137[2:2];
    assign _1412 = _137[1:1];
    assign _1411 = _137[0:0];
    assign _1423 = { _1411, _1412, _1413, _1414, _1415, _1416, _1417, _1418, _1419, _1420, _1421, _1422 };
    assign address_77 = PHASE_17 ? _60 : _1423;
    assign _1408 = ~ PHASE_17;
    assign read_enable_63 = _102 & _1408;
    assign _1406 = _62[1:1];
    assign write_enable_77 = _1406 & PHASE_17;
    assign _1410 = write_enable_77 | read_enable_63;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_37
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1410), .regcea(vdd), .wea(write_enable_77), .addra(address_77), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_62), .regceb(vdd), .web(write_enable_76), .addrb(address_76), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1445[131:131]), .sbiterrb(_1445[130:130]), .doutb(_1445[129:66]), .dbiterra(_1445[65:65]), .sbiterra(_1445[64:64]), .douta(_1445[63:0]) );
    assign _1446 = _1445[63:0];
    assign _1367 = ~ PHASE_17;
    assign _51 = _1367;
    always @(posedge _84) begin
        if (_82)
            PHASE_17 <= _1365;
        else
            if (_72)
                PHASE_17 <= _51;
    end
    assign _1460 = PHASE_17 ? _1459 : _1446;
    assign address_78 = _1391 ? _199 : _172;
    assign _1398 = ~ _1391;
    assign read_enable_64 = _102 & _1398;
    assign write_enable_78 = _1382 & _1391;
    assign _1400 = write_enable_78 | read_enable_64;
    assign address_79 = _1391 ? _164 : _137;
    assign _1393 = ~ _1391;
    assign read_enable_65 = _102 & _1393;
    assign _1391 = ~ PHASE_18;
    assign write_enable_79 = _1375 & _1391;
    assign _1395 = write_enable_79 | read_enable_65;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_38
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1395), .regcea(vdd), .wea(write_enable_79), .addra(address_79), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1400), .regceb(vdd), .web(write_enable_78), .addrb(address_78), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1403[131:131]), .sbiterrb(_1403[130:130]), .doutb(_1403[129:66]), .dbiterra(_1403[65:65]), .sbiterra(_1403[64:64]), .douta(_1403[63:0]) );
    assign _1404 = _1403[63:0];
    assign _1471 = _1470[127:64];
    assign data_75 = _1471;
    assign address_80 = PHASE_18 ? _199 : _172;
    assign _1384 = ~ PHASE_18;
    assign read_enable_66 = _102 & _1384;
    assign _1381 = ~ _130;
    assign _1382 = _129 & _1381;
    assign write_enable_80 = _1382 & PHASE_18;
    assign _1386 = write_enable_80 | read_enable_66;
    assign address_81 = PHASE_18 ? _164 : _137;
    assign _1377 = ~ PHASE_18;
    assign read_enable_67 = _102 & _1377;
    assign _1374 = ~ _130;
    assign _1375 = _129 & _1374;
    assign write_enable_81 = _1375 & PHASE_18;
    assign _1379 = write_enable_81 | read_enable_67;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_39
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1379), .regcea(vdd), .wea(write_enable_81), .addra(address_81), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1386), .regceb(vdd), .web(write_enable_80), .addrb(address_80), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1389[131:131]), .sbiterrb(_1389[130:130]), .doutb(_1389[129:66]), .dbiterra(_1389[65:65]), .sbiterra(_1389[64:64]), .douta(_1389[63:0]) );
    assign _1390 = _1389[63:0];
    assign _1472 = ~ PHASE_18;
    assign _53 = _1472;
    always @(posedge _84) begin
        if (_82)
            PHASE_18 <= _1372;
        else
            if (_99)
                PHASE_18 <= _53;
    end
    assign q0_5 = PHASE_18 ? _1404 : _1390;
    always @(posedge _84) begin
        if (_82)
            _1370 <= _1369;
        else
            _1370 <= _92;
    end
    assign _1461 = _1370 ? _1460 : q0_5;
    dp_48
        dp_0
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1461), .d2(_1468), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1470[191:128]), .q2(_1470[127:64]), .q1(_1470[63:0]) );
    assign _1473 = _1470[63:0];
    assign data_79 = _1473;
    assign address_82 = PHASE_19 ? _164 : _68;
    assign _1537 = ~ PHASE_19;
    assign _1536 = _70[1:1];
    assign read_enable_68 = _1536 & _1537;
    always @(posedge _84) begin
        if (_82)
            _1507 <= _1506;
        else
            _1507 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1510 <= _1509;
        else
            _1510 <= _1507;
    end
    always @(posedge _84) begin
        if (_82)
            _1513 <= _1512;
        else
            _1513 <= _1510;
    end
    always @(posedge _84) begin
        if (_82)
            _1516 <= _1515;
        else
            _1516 <= _1513;
    end
    always @(posedge _84) begin
        if (_82)
            _1519 <= _1518;
        else
            _1519 <= _1516;
    end
    always @(posedge _84) begin
        if (_82)
            _1522 <= _1521;
        else
            _1522 <= _1519;
    end
    always @(posedge _84) begin
        if (_82)
            _1525 <= _1524;
        else
            _1525 <= _1522;
    end
    always @(posedge _84) begin
        if (_82)
            _1528 <= _1527;
        else
            _1528 <= _1525;
    end
    always @(posedge _84) begin
        if (_82)
            _1531 <= _1530;
        else
            _1531 <= _1528;
    end
    assign _1532 = ~ _1531;
    always @(posedge _84) begin
        if (_82)
            _1480 <= _1479;
        else
            _1480 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1483 <= _1482;
        else
            _1483 <= _1480;
    end
    always @(posedge _84) begin
        if (_82)
            _1486 <= _1485;
        else
            _1486 <= _1483;
    end
    always @(posedge _84) begin
        if (_82)
            _1489 <= _1488;
        else
            _1489 <= _1486;
    end
    always @(posedge _84) begin
        if (_82)
            _1492 <= _1491;
        else
            _1492 <= _1489;
    end
    always @(posedge _84) begin
        if (_82)
            _1495 <= _1494;
        else
            _1495 <= _1492;
    end
    always @(posedge _84) begin
        if (_82)
            _1498 <= _1497;
        else
            _1498 <= _1495;
    end
    always @(posedge _84) begin
        if (_82)
            _1501 <= _1500;
        else
            _1501 <= _1498;
    end
    always @(posedge _84) begin
        if (_82)
            _1504 <= _1503;
        else
            _1504 <= _1501;
    end
    assign _1533 = _1504 & _1532;
    assign _1534 = _129 & _1533;
    assign write_enable_82 = _1534 & PHASE_19;
    assign _1539 = write_enable_82 | read_enable_68;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_40
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1539), .regcea(vdd), .wea(write_enable_82), .addra(address_82), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_73), .regceb(vdd), .web(write_enable_73), .addrb(address_73), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1546[131:131]), .sbiterrb(_1546[130:130]), .doutb(_1546[129:66]), .dbiterra(_1546[65:65]), .sbiterra(_1546[64:64]), .douta(_1546[63:0]) );
    assign _1547 = _1546[63:0];
    assign _1477 = ~ PHASE_19;
    assign _55 = _1477;
    always @(posedge _84) begin
        if (_82)
            PHASE_19 <= _1475;
        else
            if (_72)
                PHASE_19 <= _55;
    end
    assign _1559 = PHASE_19 ? _1558 : _1547;
    assign address_83 = _1744 ? _199 : _1739;
    assign write_enable_83 = _1737 & _1744;
    assign address_84 = _1744 ? _164 : _68;
    assign _1746 = ~ _1744;
    assign read_enable_69 = _1732 & _1746;
    assign _1744 = ~ PHASE_22;
    assign write_enable_84 = _1730 & _1744;
    assign _1748 = write_enable_84 | read_enable_69;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_41
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1748), .regcea(vdd), .wea(write_enable_84), .addra(address_84), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_83), .regceb(vdd), .web(write_enable_83), .addrb(address_83), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1753[131:131]), .sbiterrb(_1753[130:130]), .doutb(_1753[129:66]), .dbiterra(_1753[65:65]), .sbiterra(_1753[64:64]), .douta(_1753[63:0]) );
    assign _1754 = _1753[63:0];
    assign address_85 = PHASE_22 ? _199 : _1739;
    assign _1737 = _129 & _1700;
    assign write_enable_85 = _1737 & PHASE_22;
    assign _292 = _91[521:518];
    assign _291 = _91[517:517];
    assign _289 = _91[513:513];
    assign _288 = _91[512:449];
    assign _287 = _91[448:385];
    assign _286 = _91[384:321];
    assign _285 = _91[320:257];
    assign _284 = _91[256:193];
    assign _283 = _91[192:129];
    assign _282 = _91[128:65];
    assign _1662 = _1654[129:66];
    assign _1661 = _1641[129:66];
    assign _1663 = PHASE_20 ? _1662 : _1661;
    assign _1659 = _1599[129:66];
    assign _1658 = _1585[129:66];
    assign q1_6 = PHASE_21 ? _1659 : _1658;
    assign _1664 = _1566 ? _1663 : q1_6;
    assign address_86 = _1643 ? _1637 : _1636;
    assign _1649 = ~ _1643;
    assign read_enable_70 = _102 & _1649;
    assign address_87 = _1643 ? _60 : _1619;
    assign _1645 = ~ _1643;
    assign read_enable_71 = _102 & _1645;
    assign _1643 = ~ PHASE_20;
    assign write_enable_87 = _1602 & _1643;
    assign _1647 = write_enable_87 | read_enable_71;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_42
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1647), .regcea(vdd), .wea(write_enable_87), .addra(address_87), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_70), .regceb(vdd), .web(write_enable_86), .addrb(address_86), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1654[131:131]), .sbiterrb(_1654[130:130]), .doutb(_1654[129:66]), .dbiterra(_1654[65:65]), .sbiterra(_1654[64:64]), .douta(_1654[63:0]) );
    assign _1655 = _1654[63:0];
    assign _1635 = _172[11:11];
    assign _1634 = _172[10:10];
    assign _1633 = _172[9:9];
    assign _1632 = _172[8:8];
    assign _1631 = _172[7:7];
    assign _1630 = _172[6:6];
    assign _1629 = _172[5:5];
    assign _1628 = _172[4:4];
    assign _1627 = _172[3:3];
    assign _1626 = _172[2:2];
    assign _1625 = _172[1:1];
    assign _1624 = _172[0:0];
    assign _1636 = { _1624, _1625, _1626, _1627, _1628, _1629, _1630, _1631, _1632, _1633, _1634, _1635 };
    assign address_88 = PHASE_20 ? _1637 : _1636;
    assign _1621 = ~ PHASE_20;
    assign read_enable_72 = _102 & _1621;
    assign data_85 = wr_d0;
    assign _60 = wr_addr;
    assign _1618 = _137[11:11];
    assign _1617 = _137[10:10];
    assign _1616 = _137[9:9];
    assign _1615 = _137[8:8];
    assign _1614 = _137[7:7];
    assign _1613 = _137[6:6];
    assign _1612 = _137[5:5];
    assign _1611 = _137[4:4];
    assign _1610 = _137[3:3];
    assign _1609 = _137[2:2];
    assign _1608 = _137[1:1];
    assign _1607 = _137[0:0];
    assign _1619 = { _1607, _1608, _1609, _1610, _1611, _1612, _1613, _1614, _1615, _1616, _1617, _1618 };
    assign address_89 = PHASE_20 ? _60 : _1619;
    assign _1604 = ~ PHASE_20;
    assign read_enable_73 = _102 & _1604;
    assign _62 = wr_en;
    assign _1602 = _62[0:0];
    assign write_enable_89 = _1602 & PHASE_20;
    assign _1606 = write_enable_89 | read_enable_73;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_43
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1606), .regcea(vdd), .wea(write_enable_89), .addra(address_89), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_72), .regceb(vdd), .web(write_enable_88), .addrb(address_88), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1641[131:131]), .sbiterrb(_1641[130:130]), .doutb(_1641[129:66]), .dbiterra(_1641[65:65]), .sbiterra(_1641[64:64]), .douta(_1641[63:0]) );
    assign _1642 = _1641[63:0];
    assign _1563 = ~ PHASE_20;
    assign _63 = _1563;
    always @(posedge _84) begin
        if (_82)
            PHASE_20 <= _1561;
        else
            if (_72)
                PHASE_20 <= _63;
    end
    assign _1656 = PHASE_20 ? _1655 : _1642;
    assign address_90 = _1587 ? _199 : _172;
    assign _1594 = ~ _1587;
    assign read_enable_74 = _102 & _1594;
    assign write_enable_90 = _1578 & _1587;
    assign _1596 = write_enable_90 | read_enable_74;
    assign address_91 = _1587 ? _164 : _137;
    assign _1589 = ~ _1587;
    assign read_enable_75 = _102 & _1589;
    assign _1587 = ~ PHASE_21;
    assign write_enable_91 = _1571 & _1587;
    assign _1591 = write_enable_91 | read_enable_75;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_44
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1591), .regcea(vdd), .wea(write_enable_91), .addra(address_91), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1596), .regceb(vdd), .web(write_enable_90), .addrb(address_90), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1599[131:131]), .sbiterrb(_1599[130:130]), .doutb(_1599[129:66]), .dbiterra(_1599[65:65]), .sbiterra(_1599[64:64]), .douta(_1599[63:0]) );
    assign _1600 = _1599[63:0];
    assign _1667 = _1666[127:64];
    assign data_87 = _1667;
    always @(posedge _84) begin
        if (_82)
            _175 <= _174;
        else
            _175 <= _172;
    end
    always @(posedge _84) begin
        if (_82)
            _178 <= _177;
        else
            _178 <= _175;
    end
    always @(posedge _84) begin
        if (_82)
            _181 <= _180;
        else
            _181 <= _178;
    end
    always @(posedge _84) begin
        if (_82)
            _184 <= _183;
        else
            _184 <= _181;
    end
    always @(posedge _84) begin
        if (_82)
            _187 <= _186;
        else
            _187 <= _184;
    end
    always @(posedge _84) begin
        if (_82)
            _190 <= _189;
        else
            _190 <= _187;
    end
    always @(posedge _84) begin
        if (_82)
            _193 <= _192;
        else
            _193 <= _190;
    end
    always @(posedge _84) begin
        if (_82)
            _196 <= _195;
        else
            _196 <= _193;
    end
    always @(posedge _84) begin
        if (_82)
            _199 <= _198;
        else
            _199 <= _196;
    end
    assign _172 = _91[64:53];
    assign address_92 = PHASE_21 ? _199 : _172;
    assign _1580 = ~ PHASE_21;
    assign read_enable_76 = _102 & _1580;
    assign _1577 = ~ _130;
    assign _1578 = _129 & _1577;
    assign write_enable_92 = _1578 & PHASE_21;
    assign _1582 = write_enable_92 | read_enable_76;
    assign address_93 = PHASE_21 ? _164 : _137;
    assign _1573 = ~ PHASE_21;
    assign read_enable_77 = _102 & _1573;
    assign _1570 = ~ _130;
    assign _1571 = _129 & _1570;
    assign write_enable_93 = _1571 & PHASE_21;
    assign _1575 = write_enable_93 | read_enable_77;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_45
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1575), .regcea(vdd), .wea(write_enable_93), .addra(address_93), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1582), .regceb(vdd), .web(write_enable_92), .addrb(address_92), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1585[131:131]), .sbiterrb(_1585[130:130]), .doutb(_1585[129:66]), .dbiterra(_1585[65:65]), .sbiterra(_1585[64:64]), .douta(_1585[63:0]) );
    assign _1586 = _1585[63:0];
    assign _99 = _91[523:523];
    assign _1668 = ~ PHASE_21;
    assign _65 = _1668;
    always @(posedge _84) begin
        if (_82)
            PHASE_21 <= _1568;
        else
            if (_99)
                PHASE_21 <= _65;
    end
    assign q0_6 = PHASE_21 ? _1600 : _1586;
    assign _92 = _91[514:514];
    always @(posedge _84) begin
        if (_82)
            _1566 <= _1565;
        else
            _1566 <= _92;
    end
    assign _1657 = _1566 ? _1656 : q0_6;
    dp_47
        dp
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1657), .d2(_1664), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1666[191:128]), .q2(_1666[127:64]), .q1(_1666[63:0]) );
    assign _1669 = _1666[63:0];
    assign data_91 = _1669;
    assign _137 = _91[52:41];
    always @(posedge _84) begin
        if (_82)
            _140 <= _139;
        else
            _140 <= _137;
    end
    always @(posedge _84) begin
        if (_82)
            _143 <= _142;
        else
            _143 <= _140;
    end
    always @(posedge _84) begin
        if (_82)
            _146 <= _145;
        else
            _146 <= _143;
    end
    always @(posedge _84) begin
        if (_82)
            _149 <= _148;
        else
            _149 <= _146;
    end
    always @(posedge _84) begin
        if (_82)
            _152 <= _151;
        else
            _152 <= _149;
    end
    always @(posedge _84) begin
        if (_82)
            _155 <= _154;
        else
            _155 <= _152;
    end
    always @(posedge _84) begin
        if (_82)
            _158 <= _157;
        else
            _158 <= _155;
    end
    always @(posedge _84) begin
        if (_82)
            _161 <= _160;
        else
            _161 <= _158;
    end
    always @(posedge _84) begin
        if (_82)
            _164 <= _163;
        else
            _164 <= _161;
    end
    assign _68 = rd_addr;
    assign address_94 = PHASE_22 ? _164 : _68;
    assign _1733 = ~ PHASE_22;
    assign _70 = rd_en;
    assign _1732 = _70[0:0];
    assign read_enable_78 = _1732 & _1733;
    assign _290 = _91[516:516];
    always @(posedge _84) begin
        if (_82)
            _1703 <= _1702;
        else
            _1703 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1706 <= _1705;
        else
            _1706 <= _1703;
    end
    always @(posedge _84) begin
        if (_82)
            _1709 <= _1708;
        else
            _1709 <= _1706;
    end
    always @(posedge _84) begin
        if (_82)
            _1712 <= _1711;
        else
            _1712 <= _1709;
    end
    always @(posedge _84) begin
        if (_82)
            _1715 <= _1714;
        else
            _1715 <= _1712;
    end
    always @(posedge _84) begin
        if (_82)
            _1718 <= _1717;
        else
            _1718 <= _1715;
    end
    always @(posedge _84) begin
        if (_82)
            _1721 <= _1720;
        else
            _1721 <= _1718;
    end
    always @(posedge _84) begin
        if (_82)
            _1724 <= _1723;
        else
            _1724 <= _1721;
    end
    always @(posedge _84) begin
        if (_82)
            _1727 <= _1726;
        else
            _1727 <= _1724;
    end
    assign _1728 = ~ _1727;
    assign _130 = _91[515:515];
    always @(posedge _84) begin
        if (_82)
            _1676 <= _1675;
        else
            _1676 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1679 <= _1678;
        else
            _1679 <= _1676;
    end
    always @(posedge _84) begin
        if (_82)
            _1682 <= _1681;
        else
            _1682 <= _1679;
    end
    always @(posedge _84) begin
        if (_82)
            _1685 <= _1684;
        else
            _1685 <= _1682;
    end
    always @(posedge _84) begin
        if (_82)
            _1688 <= _1687;
        else
            _1688 <= _1685;
    end
    always @(posedge _84) begin
        if (_82)
            _1691 <= _1690;
        else
            _1691 <= _1688;
    end
    always @(posedge _84) begin
        if (_82)
            _1694 <= _1693;
        else
            _1694 <= _1691;
    end
    always @(posedge _84) begin
        if (_82)
            _1697 <= _1696;
        else
            _1697 <= _1694;
    end
    always @(posedge _84) begin
        if (_82)
            _1700 <= _1699;
        else
            _1700 <= _1697;
    end
    assign _1729 = _1700 & _1728;
    assign _102 = _91[522:522];
    always @(posedge _84) begin
        if (_82)
            _105 <= _104;
        else
            _105 <= _102;
    end
    always @(posedge _84) begin
        if (_82)
            _108 <= _107;
        else
            _108 <= _105;
    end
    always @(posedge _84) begin
        if (_82)
            _111 <= _110;
        else
            _111 <= _108;
    end
    always @(posedge _84) begin
        if (_82)
            _114 <= _113;
        else
            _114 <= _111;
    end
    always @(posedge _84) begin
        if (_82)
            _117 <= _116;
        else
            _117 <= _114;
    end
    always @(posedge _84) begin
        if (_82)
            _120 <= _119;
        else
            _120 <= _117;
    end
    always @(posedge _84) begin
        if (_82)
            _123 <= _122;
        else
            _123 <= _120;
    end
    always @(posedge _84) begin
        if (_82)
            _126 <= _125;
        else
            _126 <= _123;
    end
    always @(posedge _84) begin
        if (_82)
            _129 <= _128;
        else
            _129 <= _126;
    end
    assign _1730 = _129 & _1729;
    assign write_enable_94 = _1730 & PHASE_22;
    assign _1735 = write_enable_94 | read_enable_78;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_46
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1735), .regcea(vdd), .wea(write_enable_94), .addra(address_94), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_85), .regceb(vdd), .web(write_enable_85), .addrb(address_85), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1742[131:131]), .sbiterrb(_1742[130:130]), .doutb(_1742[129:66]), .dbiterra(_1742[65:65]), .sbiterra(_1742[64:64]), .douta(_1742[63:0]) );
    assign _1743 = _1742[63:0];
    assign _72 = flip;
    assign _1673 = ~ PHASE_22;
    assign _73 = _1673;
    always @(posedge _84) begin
        if (_82)
            PHASE_22 <= _1671;
        else
            if (_72)
                PHASE_22 <= _73;
    end
    assign _1755 = PHASE_22 ? _1754 : _1743;
    assign _76 = first_4step_pass;
    assign _78 = first_iter;
    assign _80 = start;
    assign _82 = clear;
    assign _84 = clock;
    ctrl
        ctrl
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .first_4step_pass(_76), .flip(_91[523:523]), .read_write_enable(_91[522:522]), .index(_91[521:518]), .valid(_91[517:517]), .twiddle_stage(_91[516:516]), .last_stage(_91[515:515]), .first_stage(_91[514:514]), .start_twiddles(_91[513:513]), .omegas6(_91[512:449]), .omegas5(_91[448:385]), .omegas4(_91[384:321]), .omegas3(_91[320:257]), .omegas2(_91[256:193]), .omegas1(_91[192:129]), .omegas0(_91[128:65]), .addr2(_91[64:53]), .addr1(_91[52:41]), .m(_91[40:29]), .k(_91[28:17]), .j(_91[16:5]), .i(_91[4:1]), .done_(_91[0:0]) );
    assign _1756 = _91[0:0];

    /* aliases */
    assign data_0 = data;
    assign data_2 = data_1;
    assign data_4 = data_3;
    assign data_5 = data_3;
    assign data_6 = data_3;
    assign data_8 = data_7;
    assign data_9 = data_7;
    assign data_10 = data_7;
    assign data_12 = data_11;
    assign data_14 = data_13;
    assign data_16 = data_15;
    assign data_17 = data_15;
    assign data_18 = data_15;
    assign data_20 = data_19;
    assign data_21 = data_19;
    assign data_22 = data_19;
    assign data_24 = data_23;
    assign data_26 = data_25;
    assign data_28 = data_27;
    assign data_29 = data_27;
    assign data_30 = data_27;
    assign data_32 = data_31;
    assign data_33 = data_31;
    assign data_34 = data_31;
    assign data_36 = data_35;
    assign data_38 = data_37;
    assign data_40 = data_39;
    assign data_41 = data_39;
    assign data_42 = data_39;
    assign data_44 = data_43;
    assign data_45 = data_43;
    assign data_46 = data_43;
    assign data_48 = data_47;
    assign data_50 = data_49;
    assign data_52 = data_51;
    assign data_53 = data_51;
    assign data_54 = data_51;
    assign data_56 = data_55;
    assign data_57 = data_55;
    assign data_58 = data_55;
    assign data_60 = data_59;
    assign data_62 = data_61;
    assign data_64 = data_63;
    assign data_65 = data_63;
    assign data_66 = data_63;
    assign data_68 = data_67;
    assign data_69 = data_67;
    assign data_70 = data_67;
    assign data_72 = data_71;
    assign data_74 = data_73;
    assign data_76 = data_75;
    assign data_77 = data_75;
    assign data_78 = data_75;
    assign data_80 = data_79;
    assign data_81 = data_79;
    assign data_82 = data_79;
    assign data_84 = data_83;
    assign data_86 = data_85;
    assign data_88 = data_87;
    assign data_89 = data_87;
    assign data_90 = data_87;
    assign data_92 = data_91;
    assign data_93 = data_91;
    assign data_94 = data_91;

    /* output assignments */
    assign done_ = _1756;
    assign rd_q0 = _1755;
    assign rd_q1 = _1559;
    assign rd_q2 = _1363;
    assign rd_q3 = _1167;
    assign rd_q4 = _971;
    assign rd_q5 = _775;
    assign rd_q6 = _579;
    assign rd_q7 = _383;

endmodule
module dp_55 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1011101011001111100011010010101101011001010000110011010011011010;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1011110000101000110110001111100101001011011110101100100100000000;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1010011101011010110000101010010100001010011101010010100011111111;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0111100010011001111011110010110000010101011010110010100000110001;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1011011110011011001100001001011100001010101001010000110000111110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0001011010011001110010100011110011001100000000011000111101010101;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0100000001000101111010011110100001010111011001101011110100011101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_56 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0001100011110101110101100101000001110101001000111100010111110100;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0011100000001010100000101010000100011110001011111111100110100001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0101011100101011100000011011010110001011100111101011010111001100;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0111001111011001100001101101101110110111101001010001010011001101;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1111001010110010100010111100011011000111001101101101110111110000;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1100100010110010000000011011001100000010111000101000000110010110;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1000101010000001010100111101100011011111111101101100100000001101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_57 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1100001111100010110101001101001100100000110100010011110110100010;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1000011011011101000110000111110111011011001000001100111111011110;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0111000111011101111101100001001011111110000010010101110010000011;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0111101101101110001011000011001010110100111001101001101110101101;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0000100110010111110010100100111100001101011111100110010000100111;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1110011011001110001111101000111100010010100010010100000110001111;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0111011001011011100010101110000100110011001100001000011000011111;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_58 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0011001000000011001110011001000010101000100000110011101101100000;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1011011011010101011100011010101010101001101001011011010100001100;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0101100100110101001011011101001001001111011001100001011101101111;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0000000111101110001110010101000001001010011000111101101011011101;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0000100100101010110101110011001010101011001010110101100100110001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0100101011001000110110011001101101111001000111110011010001101001;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0010110100011001110001010100101100111100010101001001010011001101;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_59 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0010100001000111001111010110011010101101010010000011001000111110;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0100010000101110000010110010110001110101010010101100101000101100;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0110011000111100001011010000011010111111001001111000111011100101;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0000010100000011100011000110011101011000001110100111010001011001;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1010101100000000110010110011010110110001111111010100000010011110;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0101001110010000111001101101001110111101111110001100111010111111;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0101100000001101011100101110110101101100101000101100101011001111;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_60 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0010100111010110111100111101011110000100010111101101111110010110;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1010010010100101001010000101110010001100011001001101101000110101;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1100000011111100110100011100010010110001000000011010010001100011;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0011010000010011111001101100101100010100011011010010001011010101;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1000011101101001011011111001101100101110001111001001110110011001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b0110011000111100000101000111101011100000110000000010010111010100;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0001100011110011100000001101000111101110001011000100011000111010;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_61 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b1111010011100010011100110010000001111101011110111111110110111011;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b1011000011111010001100001001100000100110100100111110101000001101;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b0010011001011100000110001010101011011111011000000001111101111000;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0011111100110001110100011101110101111111111110110000010011010110;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b0011000010001100001100011100100111111111000000110100110000111001;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1001000110010011001111101000110110101010110010001101001001001111;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b1101101111001011010111001011111000101000101010100101110101010110;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module dp_62 (
    omegas6,
    omegas5,
    omegas4,
    omegas3,
    omegas2,
    omegas1,
    omegas0,
    twiddle_stage,
    start_twiddles,
    first_iter,
    start,
    clear,
    index,
    d2,
    valid,
    clock,
    d1,
    q1,
    q2,
    twiddle_update_q
);

    input [63:0] omegas6;
    input [63:0] omegas5;
    input [63:0] omegas4;
    input [63:0] omegas3;
    input [63:0] omegas2;
    input [63:0] omegas1;
    input [63:0] omegas0;
    input twiddle_stage;
    input start_twiddles;
    input first_iter;
    input start;
    input clear;
    input [3:0] index;
    input [63:0] d2;
    input valid;
    input clock;
    input [63:0] d1;
    output [63:0] q1;
    output [63:0] q2;
    output [63:0] twiddle_update_q;

    /* signal declarations */
    wire [63:0] _104 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _103 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _98 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _99;
    wire [64:0] _95;
    wire [64:0] _94;
    wire [64:0] _96;
    wire _97;
    wire [64:0] _100;
    wire [63:0] _101;
    wire _70 = 1'b0;
    wire _69 = 1'b0;
    wire _67 = 1'b0;
    wire _66 = 1'b0;
    wire _64 = 1'b0;
    wire _63 = 1'b0;
    wire _61 = 1'b0;
    wire _60 = 1'b0;
    wire _58 = 1'b0;
    wire _57 = 1'b0;
    wire _55 = 1'b0;
    wire _54 = 1'b0;
    wire _52 = 1'b0;
    wire _51 = 1'b0;
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    reg _50;
    reg _53;
    reg _56;
    reg _59;
    reg _62;
    reg _65;
    reg _68;
    reg piped_twiddle_stage;
    wire [63:0] _102;
    reg [63:0] _105;
    wire [63:0] _295 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _294 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _290 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _291;
    wire [64:0] _287 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [63:0] _282 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _281 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _277 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _278;
    wire [64:0] _274 = 65'b01111111111111111111111111111111100000000000000000000000000000001;
    wire [64:0] _271 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _270 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [32:0] _267 = 33'b000000000000000000000000000000000;
    wire [64:0] _268;
    wire [31:0] _264 = 32'b00000000000000000000000000000000;
    wire [31:0] _263;
    wire [63:0] _265;
    wire [64:0] _266;
    wire [64:0] _269;
    reg [64:0] _272;
    wire [64:0] _261 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _260 = 65'b00000000000000000000000000000000000000000000000000000000000000000;
    wire [64:0] _257 = 65'b00000000000000000000000000000000011111111111111111111111111111111;
    wire [63:0] _255;
    wire [64:0] _256;
    wire [64:0] _258;
    wire [31:0] _251;
    wire [32:0] _250 = 33'b000000000000000000000000000000000;
    wire [64:0] _252;
    wire [127:0] _246 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _245 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _243 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _242 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _240 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [127:0] _239 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _236 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _232 = 64'b1000010001110111011101111010001101011010001110110100010100111111;
    wire [63:0] _231 = 64'b1010011111111000011110110001100010101001010001001001111110101011;
    wire [63:0] _230 = 64'b1011000000010011100110100001111101100101110000111000010011000111;
    wire [63:0] _229 = 64'b0101010011011111100101100011000010111111011110010100010100001110;
    wire [63:0] _228 = 64'b1110111111010010011111010110001000110000011000111111011001111110;
    wire [63:0] _227 = 64'b1010101111010000101001101110100010101010001111011000101000001110;
    wire [63:0] _226 = 64'b1000000100101000000110100111101100000101111110011011111010101100;
    reg [63:0] twiddle_scale;
    wire [63:0] _4;
    wire _152 = 1'b0;
    wire _151 = 1'b0;
    reg _153;
    wire [63:0] _157;
    wire [63:0] _6;
    wire _145 = 1'b0;
    wire _144 = 1'b0;
    reg _146;
    wire [63:0] _150;
    wire [63:0] _8;
    wire _138 = 1'b0;
    wire _137 = 1'b0;
    reg _139;
    wire [63:0] _143;
    wire [63:0] _10;
    wire _131 = 1'b0;
    wire _130 = 1'b0;
    reg _132;
    wire [63:0] _136;
    wire [63:0] _12;
    wire _124 = 1'b0;
    wire _123 = 1'b0;
    reg _125;
    wire [63:0] _129;
    wire [63:0] _14;
    wire _117 = 1'b0;
    wire _116 = 1'b0;
    reg _118;
    wire [63:0] _122;
    wire [63:0] _16;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _18;
    reg _111;
    wire [63:0] _115;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire _20;
    reg _108;
    wire [63:0] _159;
    wire [63:0] w;
    wire [63:0] twiddle_factor;
    wire [63:0] b;
    reg [63:0] _237;
    wire [63:0] _224 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _223 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _113 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _112 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _120 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _119 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _127 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _126 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _134 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _133 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _141 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _140 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _148 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _147 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _155 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _154 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _185 = 64'b0101000011110101101000010110011100001110011110100110000110000000;
    wire [63:0] _186;
    wire [63:0] _187;
    wire [63:0] _22;
    reg [63:0] twiddle_omega6;
    wire [63:0] _188 = 64'b0011011011110011000011111101110100101011011111110100100011001001;
    wire [63:0] _189;
    wire [63:0] _190;
    wire [63:0] _23;
    reg [63:0] twiddle_omega5;
    wire [63:0] _191 = 64'b1100101001000111101011100101000000010101001011001001001000010000;
    wire [63:0] _192;
    wire [63:0] _193;
    wire [63:0] _24;
    reg [63:0] twiddle_omega4;
    wire [63:0] _194 = 64'b0011000101111100111000111101000110001100011110101101101000010101;
    wire [63:0] _195;
    wire [63:0] _196;
    wire [63:0] _25;
    reg [63:0] twiddle_omega3;
    wire [63:0] _197 = 64'b1000110100110000010001100011010110011011111001000111010101101011;
    wire [63:0] _198;
    wire [63:0] _199;
    wire [63:0] _26;
    reg [63:0] twiddle_omega2;
    wire [63:0] _200 = 64'b1110000101110100011000000100000100110100000010000010100100010011;
    wire [63:0] _201;
    wire [63:0] _202;
    wire [63:0] _27;
    reg [63:0] twiddle_omega1;
    wire [63:0] _203 = 64'b0000010100100101000010101011110010110110000000011111001101101000;
    wire _29;
    wire _31;
    wire _184;
    wire [63:0] _204;
    wire _182 = 1'b0;
    wire _181 = 1'b0;
    wire _179 = 1'b0;
    wire _178 = 1'b0;
    wire _176 = 1'b0;
    wire _175 = 1'b0;
    wire _173 = 1'b0;
    wire _172 = 1'b0;
    wire _170 = 1'b0;
    wire _169 = 1'b0;
    wire _167 = 1'b0;
    wire _166 = 1'b0;
    wire _164 = 1'b0;
    wire _163 = 1'b0;
    wire _161 = 1'b0;
    wire _33;
    wire _160 = 1'b0;
    reg _162;
    reg _165;
    reg _168;
    reg _171;
    reg _174;
    reg _177;
    reg _180;
    reg _183;
    wire [63:0] _205;
    wire [63:0] _34;
    reg [63:0] twiddle_omega0;
    wire [3:0] _219 = 4'b0000;
    wire [3:0] _218 = 4'b0000;
    wire [3:0] _216 = 4'b0000;
    wire [3:0] _215 = 4'b0000;
    wire [3:0] _36;
    reg [3:0] _217;
    reg [3:0] _220;
    reg [63:0] _221;
    wire [63:0] _213 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _212 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _38;
    reg [63:0] piped_d2;
    wire _210 = 1'b0;
    wire _209 = 1'b0;
    wire _207 = 1'b0;
    wire _206 = 1'b0;
    wire _40;
    reg _208;
    reg piped_twidle_updated_valid;
    wire [63:0] a;
    reg [63:0] _225;
    wire [127:0] _238;
    reg [127:0] _241;
    reg [127:0] _244;
    reg [127:0] _247;
    wire [63:0] _248;
    wire [64:0] _249;
    wire [64:0] _253;
    wire _254;
    wire [64:0] _259;
    reg [64:0] _262;
    wire [64:0] _273;
    wire _275;
    wire _276;
    wire [64:0] _279;
    wire [63:0] _280;
    reg [63:0] _283;
    wire [63:0] T;
    wire [64:0] _285;
    wire [63:0] _92 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _91 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _89 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _88 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _86 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _85 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _82 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _80 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _79 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _77 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _76 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [63:0] _74 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _73 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire _43;
    wire [63:0] _45;
    reg [63:0] _75;
    reg [63:0] _78;
    reg [63:0] _81;
    reg [63:0] _84;
    reg [63:0] _87;
    reg [63:0] _90;
    reg [63:0] _93;
    wire gnd = 1'b0;
    wire [64:0] _284;
    wire [64:0] _286;
    wire _288;
    wire _289;
    wire [64:0] _292;
    wire [63:0] _293;
    reg [63:0] _296;

    /* logic */
    assign _99 = _96 + _98;
    assign _95 = { gnd, T };
    assign _94 = { gnd, _93 };
    assign _96 = _94 - _95;
    assign _97 = _96[64:64];
    assign _100 = _97 ? _99 : _96;
    assign _101 = _100[63:0];
    always @(posedge _43) begin
        _50 <= _18;
    end
    always @(posedge _43) begin
        _53 <= _50;
    end
    always @(posedge _43) begin
        _56 <= _53;
    end
    always @(posedge _43) begin
        _59 <= _56;
    end
    always @(posedge _43) begin
        _62 <= _59;
    end
    always @(posedge _43) begin
        _65 <= _62;
    end
    always @(posedge _43) begin
        _68 <= _65;
    end
    always @(posedge _43) begin
        piped_twiddle_stage <= _68;
    end
    assign _102 = piped_twiddle_stage ? T : _101;
    always @(posedge _43) begin
        _105 <= _102;
    end
    assign _291 = _286 - _290;
    assign _278 = _273 - _277;
    assign _268 = { _267, _263 };
    assign _263 = _247[95:64];
    assign _265 = { _263, _264 };
    assign _266 = { gnd, _265 };
    assign _269 = _266 - _268;
    always @(posedge _43) begin
        _272 <= _269;
    end
    assign _255 = _253[63:0];
    assign _256 = { gnd, _255 };
    assign _258 = _256 - _257;
    assign _251 = _247[127:96];
    assign _252 = { _250, _251 };
    always @* begin
        case (_220)
        0: twiddle_scale <= _226;
        1: twiddle_scale <= _227;
        2: twiddle_scale <= _228;
        3: twiddle_scale <= _229;
        4: twiddle_scale <= _230;
        5: twiddle_scale <= _231;
        default: twiddle_scale <= _232;
        endcase
    end
    assign _4 = omegas6;
    always @(posedge _43) begin
        _153 <= _18;
    end
    assign _157 = _153 ? twiddle_omega6 : _4;
    assign _6 = omegas5;
    always @(posedge _43) begin
        _146 <= _18;
    end
    assign _150 = _146 ? twiddle_omega5 : _6;
    assign _8 = omegas4;
    always @(posedge _43) begin
        _139 <= _18;
    end
    assign _143 = _139 ? twiddle_omega4 : _8;
    assign _10 = omegas3;
    always @(posedge _43) begin
        _132 <= _18;
    end
    assign _136 = _132 ? twiddle_omega3 : _10;
    assign _12 = omegas2;
    always @(posedge _43) begin
        _125 <= _18;
    end
    assign _129 = _125 ? twiddle_omega2 : _12;
    assign _14 = omegas1;
    always @(posedge _43) begin
        _118 <= _18;
    end
    assign _122 = _118 ? twiddle_omega1 : _14;
    assign _16 = omegas0;
    assign _18 = twiddle_stage;
    always @(posedge _43) begin
        _111 <= _18;
    end
    assign _115 = _111 ? twiddle_omega0 : _16;
    assign _20 = start_twiddles;
    always @(posedge _43) begin
        if (_33)
            _108 <= _107;
        else
            _108 <= _20;
    end
    twdl
        twdl
        ( .clock(_43), .start_twiddles(_108), .omegas0(_115), .omegas1(_122), .omegas2(_129), .omegas3(_136), .omegas4(_143), .omegas5(_150), .omegas6(_157), .w(_159[63:0]) );
    assign w = _159;
    assign b = piped_twidle_updated_valid ? twiddle_scale : w;
    always @(posedge _43) begin
        _237 <= b;
    end
    assign _186 = _184 ? _185 : twiddle_omega6;
    assign _187 = _183 ? T : _186;
    assign _22 = _187;
    always @(posedge _43) begin
        twiddle_omega6 <= _22;
    end
    assign _189 = _184 ? _188 : twiddle_omega5;
    assign _190 = _183 ? twiddle_omega6 : _189;
    assign _23 = _190;
    always @(posedge _43) begin
        twiddle_omega5 <= _23;
    end
    assign _192 = _184 ? _191 : twiddle_omega4;
    assign _193 = _183 ? twiddle_omega5 : _192;
    assign _24 = _193;
    always @(posedge _43) begin
        twiddle_omega4 <= _24;
    end
    assign _195 = _184 ? _194 : twiddle_omega3;
    assign _196 = _183 ? twiddle_omega4 : _195;
    assign _25 = _196;
    always @(posedge _43) begin
        twiddle_omega3 <= _25;
    end
    assign _198 = _184 ? _197 : twiddle_omega2;
    assign _199 = _183 ? twiddle_omega3 : _198;
    assign _26 = _199;
    always @(posedge _43) begin
        twiddle_omega2 <= _26;
    end
    assign _201 = _184 ? _200 : twiddle_omega1;
    assign _202 = _183 ? twiddle_omega2 : _201;
    assign _27 = _202;
    always @(posedge _43) begin
        twiddle_omega1 <= _27;
    end
    assign _29 = first_iter;
    assign _31 = start;
    assign _184 = _31 & _29;
    assign _204 = _184 ? _203 : twiddle_omega0;
    assign _33 = clear;
    always @(posedge _43) begin
        if (_33)
            _162 <= _161;
        else
            _162 <= _40;
    end
    always @(posedge _43) begin
        if (_33)
            _165 <= _164;
        else
            _165 <= _162;
    end
    always @(posedge _43) begin
        if (_33)
            _168 <= _167;
        else
            _168 <= _165;
    end
    always @(posedge _43) begin
        if (_33)
            _171 <= _170;
        else
            _171 <= _168;
    end
    always @(posedge _43) begin
        if (_33)
            _174 <= _173;
        else
            _174 <= _171;
    end
    always @(posedge _43) begin
        if (_33)
            _177 <= _176;
        else
            _177 <= _174;
    end
    always @(posedge _43) begin
        if (_33)
            _180 <= _179;
        else
            _180 <= _177;
    end
    always @(posedge _43) begin
        if (_33)
            _183 <= _182;
        else
            _183 <= _180;
    end
    assign _205 = _183 ? twiddle_omega1 : _204;
    assign _34 = _205;
    always @(posedge _43) begin
        twiddle_omega0 <= _34;
    end
    assign _36 = index;
    always @(posedge _43) begin
        _217 <= _36;
    end
    always @(posedge _43) begin
        _220 <= _217;
    end
    always @* begin
        case (_220)
        0: _221 <= twiddle_omega0;
        1: _221 <= twiddle_omega1;
        2: _221 <= twiddle_omega2;
        3: _221 <= twiddle_omega3;
        4: _221 <= twiddle_omega4;
        5: _221 <= twiddle_omega5;
        default: _221 <= twiddle_omega6;
        endcase
    end
    assign _38 = d2;
    always @(posedge _43) begin
        piped_d2 <= _38;
    end
    assign _40 = valid;
    always @(posedge _43) begin
        _208 <= _40;
    end
    always @(posedge _43) begin
        piped_twidle_updated_valid <= _208;
    end
    assign a = piped_twidle_updated_valid ? _221 : piped_d2;
    always @(posedge _43) begin
        _225 <= a;
    end
    assign _238 = _225 * _237;
    always @(posedge _43) begin
        _241 <= _238;
    end
    always @(posedge _43) begin
        _244 <= _241;
    end
    always @(posedge _43) begin
        _247 <= _244;
    end
    assign _248 = _247[63:0];
    assign _249 = { gnd, _248 };
    assign _253 = _249 - _252;
    assign _254 = _253[64:64];
    assign _259 = _254 ? _258 : _253;
    always @(posedge _43) begin
        _262 <= _259;
    end
    assign _273 = _262 + _272;
    assign _275 = _273 < _274;
    assign _276 = ~ _275;
    assign _279 = _276 ? _278 : _273;
    assign _280 = _279[63:0];
    always @(posedge _43) begin
        _283 <= _280;
    end
    assign T = _283;
    assign _285 = { gnd, T };
    assign _43 = clock;
    assign _45 = d1;
    always @(posedge _43) begin
        _75 <= _45;
    end
    always @(posedge _43) begin
        _78 <= _75;
    end
    always @(posedge _43) begin
        _81 <= _78;
    end
    always @(posedge _43) begin
        _84 <= _81;
    end
    always @(posedge _43) begin
        _87 <= _84;
    end
    always @(posedge _43) begin
        _90 <= _87;
    end
    always @(posedge _43) begin
        _93 <= _90;
    end
    assign _284 = { gnd, _93 };
    assign _286 = _284 + _285;
    assign _288 = _286 < _287;
    assign _289 = ~ _288;
    assign _292 = _289 ? _291 : _286;
    assign _293 = _292[63:0];
    always @(posedge _43) begin
        _296 <= _293;
    end

    /* aliases */
    assign twiddle_factor = w;

    /* output assignments */
    assign q1 = _296;
    assign q2 = _105;
    assign twiddle_update_q = T;

endmodule
module parallel_cores_6 (
    wr_d7,
    wr_d6,
    wr_d5,
    wr_d4,
    wr_d3,
    wr_d2,
    wr_d1,
    wr_d0,
    wr_addr,
    wr_en,
    rd_addr,
    rd_en,
    flip,
    first_4step_pass,
    first_iter,
    start,
    clear,
    clock,
    done_,
    rd_q0,
    rd_q1,
    rd_q2,
    rd_q3,
    rd_q4,
    rd_q5,
    rd_q6,
    rd_q7
);

    input [63:0] wr_d7;
    input [63:0] wr_d6;
    input [63:0] wr_d5;
    input [63:0] wr_d4;
    input [63:0] wr_d3;
    input [63:0] wr_d2;
    input [63:0] wr_d1;
    input [63:0] wr_d0;
    input [11:0] wr_addr;
    input [7:0] wr_en;
    input [11:0] rd_addr;
    input [7:0] rd_en;
    input flip;
    input first_4step_pass;
    input first_iter;
    input start;
    input clear;
    input clock;
    output done_;
    output [63:0] rd_q0;
    output [63:0] rd_q1;
    output [63:0] rd_q2;
    output [63:0] rd_q3;
    output [63:0] rd_q4;
    output [63:0] rd_q5;
    output [63:0] rd_q6;
    output [63:0] rd_q7;

    /* signal declarations */
    wire [11:0] address;
    wire write_enable;
    wire [11:0] address_0;
    wire _374;
    wire read_enable;
    wire _372;
    wire write_enable_0;
    wire _376;
    wire [131:0] _381;
    wire [63:0] _382;
    wire [11:0] _367 = 12'b000000000000;
    wire [11:0] address_1;
    wire _365;
    wire write_enable_1;
    wire [63:0] _279;
    wire [63:0] _278;
    wire [63:0] _280;
    wire [63:0] _276;
    wire [63:0] _275;
    wire [63:0] q1;
    wire [63:0] _281;
    wire [11:0] address_2;
    wire write_enable_2 = 1'b0;
    wire _266;
    wire read_enable_0;
    wire [11:0] address_3;
    wire _262;
    wire read_enable_1;
    wire _260;
    wire write_enable_3;
    wire _264;
    wire [131:0] _271;
    wire [63:0] _272;
    wire [63:0] data = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_0;
    wire [11:0] _254 = 12'b000000000000;
    wire _252;
    wire _251;
    wire _250;
    wire _249;
    wire _248;
    wire _247;
    wire _246;
    wire _245;
    wire _244;
    wire _243;
    wire _242;
    wire _241;
    wire [11:0] _253;
    wire [11:0] address_4;
    wire write_enable_4 = 1'b0;
    wire _238;
    wire read_enable_2;
    wire [63:0] data_1;
    wire [63:0] data_2;
    wire _235;
    wire _234;
    wire _233;
    wire _232;
    wire _231;
    wire _230;
    wire _229;
    wire _228;
    wire _227;
    wire _226;
    wire _225;
    wire _224;
    wire [11:0] _236;
    wire [11:0] address_5;
    wire _221;
    wire read_enable_3;
    wire _219;
    wire write_enable_5;
    wire _223;
    wire [131:0] _258;
    wire [63:0] _259;
    wire _87 = 1'b0;
    wire _86 = 1'b0;
    wire _89;
    wire _3;
    reg PHASE;
    wire [63:0] _273;
    wire [11:0] address_6;
    wire _211;
    wire read_enable_4;
    wire write_enable_6;
    wire _213;
    wire [11:0] address_7;
    wire _206;
    wire read_enable_5;
    wire _204;
    wire write_enable_7;
    wire _208;
    wire [131:0] _216;
    wire [63:0] _217;
    wire [63:0] _295;
    wire [63:0] data_3;
    wire [63:0] data_4;
    wire [63:0] data_5;
    wire [63:0] data_6;
    wire [11:0] address_8;
    wire _169;
    wire read_enable_6;
    wire _166;
    wire _167;
    wire write_enable_8;
    wire _171;
    wire [11:0] address_9;
    wire _134;
    wire read_enable_7;
    wire _131;
    wire _132;
    wire write_enable_9;
    wire _136;
    wire [131:0] _202;
    wire [63:0] _203;
    wire _98 = 1'b0;
    wire _97 = 1'b0;
    wire _296;
    wire _5;
    reg PHASE_0;
    wire [63:0] q0;
    wire _94 = 1'b0;
    wire _93 = 1'b0;
    reg _96;
    wire [63:0] _274;
    wire [191:0] _294;
    wire [63:0] _297;
    wire [63:0] data_7;
    wire [63:0] data_8;
    wire [63:0] data_9;
    wire [63:0] data_10;
    wire [11:0] address_10;
    wire _361;
    wire _360;
    wire read_enable_8;
    wire _354 = 1'b0;
    wire _353 = 1'b0;
    wire _351 = 1'b0;
    wire _350 = 1'b0;
    wire _348 = 1'b0;
    wire _347 = 1'b0;
    wire _345 = 1'b0;
    wire _344 = 1'b0;
    wire _342 = 1'b0;
    wire _341 = 1'b0;
    wire _339 = 1'b0;
    wire _338 = 1'b0;
    wire _336 = 1'b0;
    wire _335 = 1'b0;
    wire _333 = 1'b0;
    wire _332 = 1'b0;
    wire _330 = 1'b0;
    wire _329 = 1'b0;
    reg _331;
    reg _334;
    reg _337;
    reg _340;
    reg _343;
    reg _346;
    reg _349;
    reg _352;
    reg _355;
    wire _356;
    wire _327 = 1'b0;
    wire _326 = 1'b0;
    wire _324 = 1'b0;
    wire _323 = 1'b0;
    wire _321 = 1'b0;
    wire _320 = 1'b0;
    wire _318 = 1'b0;
    wire _317 = 1'b0;
    wire _315 = 1'b0;
    wire _314 = 1'b0;
    wire _312 = 1'b0;
    wire _311 = 1'b0;
    wire _309 = 1'b0;
    wire _308 = 1'b0;
    wire _306 = 1'b0;
    wire _305 = 1'b0;
    wire _303 = 1'b0;
    wire _302 = 1'b0;
    reg _304;
    reg _307;
    reg _310;
    reg _313;
    reg _316;
    reg _319;
    reg _322;
    reg _325;
    reg _328;
    wire _357;
    wire _358;
    wire write_enable_10;
    wire _363;
    wire [131:0] _370;
    wire [63:0] _371;
    wire _299 = 1'b0;
    wire _298 = 1'b0;
    wire _301;
    wire _7;
    reg PHASE_1;
    wire [63:0] _383;
    wire [11:0] address_11;
    wire write_enable_11;
    wire [11:0] address_12;
    wire _570;
    wire read_enable_9;
    wire _568;
    wire write_enable_12;
    wire _572;
    wire [131:0] _577;
    wire [63:0] _578;
    wire [11:0] _563 = 12'b000000000000;
    wire [11:0] address_13;
    wire _561;
    wire write_enable_13;
    wire [63:0] _486;
    wire [63:0] _485;
    wire [63:0] _487;
    wire [63:0] _483;
    wire [63:0] _482;
    wire [63:0] q1_0;
    wire [63:0] _488;
    wire [11:0] address_14;
    wire write_enable_14 = 1'b0;
    wire _473;
    wire read_enable_10;
    wire [11:0] address_15;
    wire _469;
    wire read_enable_11;
    wire _467;
    wire write_enable_15;
    wire _471;
    wire [131:0] _478;
    wire [63:0] _479;
    wire [63:0] data_11 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_12;
    wire [11:0] _461 = 12'b000000000000;
    wire _459;
    wire _458;
    wire _457;
    wire _456;
    wire _455;
    wire _454;
    wire _453;
    wire _452;
    wire _451;
    wire _450;
    wire _449;
    wire _448;
    wire [11:0] _460;
    wire [11:0] address_16;
    wire write_enable_16 = 1'b0;
    wire _445;
    wire read_enable_12;
    wire [63:0] data_13;
    wire [63:0] data_14;
    wire _442;
    wire _441;
    wire _440;
    wire _439;
    wire _438;
    wire _437;
    wire _436;
    wire _435;
    wire _434;
    wire _433;
    wire _432;
    wire _431;
    wire [11:0] _443;
    wire [11:0] address_17;
    wire _428;
    wire read_enable_13;
    wire _426;
    wire write_enable_17;
    wire _430;
    wire [131:0] _465;
    wire [63:0] _466;
    wire _385 = 1'b0;
    wire _384 = 1'b0;
    wire _387;
    wire _11;
    reg PHASE_2;
    wire [63:0] _480;
    wire [11:0] address_18;
    wire _418;
    wire read_enable_14;
    wire write_enable_18;
    wire _420;
    wire [11:0] address_19;
    wire _413;
    wire read_enable_15;
    wire _411;
    wire write_enable_19;
    wire _415;
    wire [131:0] _423;
    wire [63:0] _424;
    wire [63:0] _491;
    wire [63:0] data_15;
    wire [63:0] data_16;
    wire [63:0] data_17;
    wire [63:0] data_18;
    wire [11:0] address_20;
    wire _404;
    wire read_enable_16;
    wire _401;
    wire _402;
    wire write_enable_20;
    wire _406;
    wire [11:0] address_21;
    wire _397;
    wire read_enable_17;
    wire _394;
    wire _395;
    wire write_enable_21;
    wire _399;
    wire [131:0] _409;
    wire [63:0] _410;
    wire _392 = 1'b0;
    wire _391 = 1'b0;
    wire _492;
    wire _13;
    reg PHASE_3;
    wire [63:0] q0_0;
    wire _389 = 1'b0;
    wire _388 = 1'b0;
    reg _390;
    wire [63:0] _481;
    wire [191:0] _490;
    wire [63:0] _493;
    wire [63:0] data_19;
    wire [63:0] data_20;
    wire [63:0] data_21;
    wire [63:0] data_22;
    wire [11:0] address_22;
    wire _557;
    wire _556;
    wire read_enable_18;
    wire _550 = 1'b0;
    wire _549 = 1'b0;
    wire _547 = 1'b0;
    wire _546 = 1'b0;
    wire _544 = 1'b0;
    wire _543 = 1'b0;
    wire _541 = 1'b0;
    wire _540 = 1'b0;
    wire _538 = 1'b0;
    wire _537 = 1'b0;
    wire _535 = 1'b0;
    wire _534 = 1'b0;
    wire _532 = 1'b0;
    wire _531 = 1'b0;
    wire _529 = 1'b0;
    wire _528 = 1'b0;
    wire _526 = 1'b0;
    wire _525 = 1'b0;
    reg _527;
    reg _530;
    reg _533;
    reg _536;
    reg _539;
    reg _542;
    reg _545;
    reg _548;
    reg _551;
    wire _552;
    wire _523 = 1'b0;
    wire _522 = 1'b0;
    wire _520 = 1'b0;
    wire _519 = 1'b0;
    wire _517 = 1'b0;
    wire _516 = 1'b0;
    wire _514 = 1'b0;
    wire _513 = 1'b0;
    wire _511 = 1'b0;
    wire _510 = 1'b0;
    wire _508 = 1'b0;
    wire _507 = 1'b0;
    wire _505 = 1'b0;
    wire _504 = 1'b0;
    wire _502 = 1'b0;
    wire _501 = 1'b0;
    wire _499 = 1'b0;
    wire _498 = 1'b0;
    reg _500;
    reg _503;
    reg _506;
    reg _509;
    reg _512;
    reg _515;
    reg _518;
    reg _521;
    reg _524;
    wire _553;
    wire _554;
    wire write_enable_22;
    wire _559;
    wire [131:0] _566;
    wire [63:0] _567;
    wire _495 = 1'b0;
    wire _494 = 1'b0;
    wire _497;
    wire _15;
    reg PHASE_4;
    wire [63:0] _579;
    wire [11:0] address_23;
    wire write_enable_23;
    wire [11:0] address_24;
    wire _766;
    wire read_enable_19;
    wire _764;
    wire write_enable_24;
    wire _768;
    wire [131:0] _773;
    wire [63:0] _774;
    wire [11:0] _759 = 12'b000000000000;
    wire [11:0] address_25;
    wire _757;
    wire write_enable_25;
    wire [63:0] _682;
    wire [63:0] _681;
    wire [63:0] _683;
    wire [63:0] _679;
    wire [63:0] _678;
    wire [63:0] q1_1;
    wire [63:0] _684;
    wire [11:0] address_26;
    wire write_enable_26 = 1'b0;
    wire _669;
    wire read_enable_20;
    wire [11:0] address_27;
    wire _665;
    wire read_enable_21;
    wire _663;
    wire write_enable_27;
    wire _667;
    wire [131:0] _674;
    wire [63:0] _675;
    wire [63:0] data_23 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_24;
    wire [11:0] _657 = 12'b000000000000;
    wire _655;
    wire _654;
    wire _653;
    wire _652;
    wire _651;
    wire _650;
    wire _649;
    wire _648;
    wire _647;
    wire _646;
    wire _645;
    wire _644;
    wire [11:0] _656;
    wire [11:0] address_28;
    wire write_enable_28 = 1'b0;
    wire _641;
    wire read_enable_22;
    wire [63:0] data_25;
    wire [63:0] data_26;
    wire _638;
    wire _637;
    wire _636;
    wire _635;
    wire _634;
    wire _633;
    wire _632;
    wire _631;
    wire _630;
    wire _629;
    wire _628;
    wire _627;
    wire [11:0] _639;
    wire [11:0] address_29;
    wire _624;
    wire read_enable_23;
    wire _622;
    wire write_enable_29;
    wire _626;
    wire [131:0] _661;
    wire [63:0] _662;
    wire _581 = 1'b0;
    wire _580 = 1'b0;
    wire _583;
    wire _19;
    reg PHASE_5;
    wire [63:0] _676;
    wire [11:0] address_30;
    wire _614;
    wire read_enable_24;
    wire write_enable_30;
    wire _616;
    wire [11:0] address_31;
    wire _609;
    wire read_enable_25;
    wire _607;
    wire write_enable_31;
    wire _611;
    wire [131:0] _619;
    wire [63:0] _620;
    wire [63:0] _687;
    wire [63:0] data_27;
    wire [63:0] data_28;
    wire [63:0] data_29;
    wire [63:0] data_30;
    wire [11:0] address_32;
    wire _600;
    wire read_enable_26;
    wire _597;
    wire _598;
    wire write_enable_32;
    wire _602;
    wire [11:0] address_33;
    wire _593;
    wire read_enable_27;
    wire _590;
    wire _591;
    wire write_enable_33;
    wire _595;
    wire [131:0] _605;
    wire [63:0] _606;
    wire _588 = 1'b0;
    wire _587 = 1'b0;
    wire _688;
    wire _21;
    reg PHASE_6;
    wire [63:0] q0_1;
    wire _585 = 1'b0;
    wire _584 = 1'b0;
    reg _586;
    wire [63:0] _677;
    wire [191:0] _686;
    wire [63:0] _689;
    wire [63:0] data_31;
    wire [63:0] data_32;
    wire [63:0] data_33;
    wire [63:0] data_34;
    wire [11:0] address_34;
    wire _753;
    wire _752;
    wire read_enable_28;
    wire _746 = 1'b0;
    wire _745 = 1'b0;
    wire _743 = 1'b0;
    wire _742 = 1'b0;
    wire _740 = 1'b0;
    wire _739 = 1'b0;
    wire _737 = 1'b0;
    wire _736 = 1'b0;
    wire _734 = 1'b0;
    wire _733 = 1'b0;
    wire _731 = 1'b0;
    wire _730 = 1'b0;
    wire _728 = 1'b0;
    wire _727 = 1'b0;
    wire _725 = 1'b0;
    wire _724 = 1'b0;
    wire _722 = 1'b0;
    wire _721 = 1'b0;
    reg _723;
    reg _726;
    reg _729;
    reg _732;
    reg _735;
    reg _738;
    reg _741;
    reg _744;
    reg _747;
    wire _748;
    wire _719 = 1'b0;
    wire _718 = 1'b0;
    wire _716 = 1'b0;
    wire _715 = 1'b0;
    wire _713 = 1'b0;
    wire _712 = 1'b0;
    wire _710 = 1'b0;
    wire _709 = 1'b0;
    wire _707 = 1'b0;
    wire _706 = 1'b0;
    wire _704 = 1'b0;
    wire _703 = 1'b0;
    wire _701 = 1'b0;
    wire _700 = 1'b0;
    wire _698 = 1'b0;
    wire _697 = 1'b0;
    wire _695 = 1'b0;
    wire _694 = 1'b0;
    reg _696;
    reg _699;
    reg _702;
    reg _705;
    reg _708;
    reg _711;
    reg _714;
    reg _717;
    reg _720;
    wire _749;
    wire _750;
    wire write_enable_34;
    wire _755;
    wire [131:0] _762;
    wire [63:0] _763;
    wire _691 = 1'b0;
    wire _690 = 1'b0;
    wire _693;
    wire _23;
    reg PHASE_7;
    wire [63:0] _775;
    wire [11:0] address_35;
    wire write_enable_35;
    wire [11:0] address_36;
    wire _962;
    wire read_enable_29;
    wire _960;
    wire write_enable_36;
    wire _964;
    wire [131:0] _969;
    wire [63:0] _970;
    wire [11:0] _955 = 12'b000000000000;
    wire [11:0] address_37;
    wire _953;
    wire write_enable_37;
    wire [63:0] _878;
    wire [63:0] _877;
    wire [63:0] _879;
    wire [63:0] _875;
    wire [63:0] _874;
    wire [63:0] q1_2;
    wire [63:0] _880;
    wire [11:0] address_38;
    wire write_enable_38 = 1'b0;
    wire _865;
    wire read_enable_30;
    wire [11:0] address_39;
    wire _861;
    wire read_enable_31;
    wire _859;
    wire write_enable_39;
    wire _863;
    wire [131:0] _870;
    wire [63:0] _871;
    wire [63:0] data_35 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_36;
    wire [11:0] _853 = 12'b000000000000;
    wire _851;
    wire _850;
    wire _849;
    wire _848;
    wire _847;
    wire _846;
    wire _845;
    wire _844;
    wire _843;
    wire _842;
    wire _841;
    wire _840;
    wire [11:0] _852;
    wire [11:0] address_40;
    wire write_enable_40 = 1'b0;
    wire _837;
    wire read_enable_32;
    wire [63:0] data_37;
    wire [63:0] data_38;
    wire _834;
    wire _833;
    wire _832;
    wire _831;
    wire _830;
    wire _829;
    wire _828;
    wire _827;
    wire _826;
    wire _825;
    wire _824;
    wire _823;
    wire [11:0] _835;
    wire [11:0] address_41;
    wire _820;
    wire read_enable_33;
    wire _818;
    wire write_enable_41;
    wire _822;
    wire [131:0] _857;
    wire [63:0] _858;
    wire _777 = 1'b0;
    wire _776 = 1'b0;
    wire _779;
    wire _27;
    reg PHASE_8;
    wire [63:0] _872;
    wire [11:0] address_42;
    wire _810;
    wire read_enable_34;
    wire write_enable_42;
    wire _812;
    wire [11:0] address_43;
    wire _805;
    wire read_enable_35;
    wire _803;
    wire write_enable_43;
    wire _807;
    wire [131:0] _815;
    wire [63:0] _816;
    wire [63:0] _883;
    wire [63:0] data_39;
    wire [63:0] data_40;
    wire [63:0] data_41;
    wire [63:0] data_42;
    wire [11:0] address_44;
    wire _796;
    wire read_enable_36;
    wire _793;
    wire _794;
    wire write_enable_44;
    wire _798;
    wire [11:0] address_45;
    wire _789;
    wire read_enable_37;
    wire _786;
    wire _787;
    wire write_enable_45;
    wire _791;
    wire [131:0] _801;
    wire [63:0] _802;
    wire _784 = 1'b0;
    wire _783 = 1'b0;
    wire _884;
    wire _29;
    reg PHASE_9;
    wire [63:0] q0_2;
    wire _781 = 1'b0;
    wire _780 = 1'b0;
    reg _782;
    wire [63:0] _873;
    wire [191:0] _882;
    wire [63:0] _885;
    wire [63:0] data_43;
    wire [63:0] data_44;
    wire [63:0] data_45;
    wire [63:0] data_46;
    wire [11:0] address_46;
    wire _949;
    wire _948;
    wire read_enable_38;
    wire _942 = 1'b0;
    wire _941 = 1'b0;
    wire _939 = 1'b0;
    wire _938 = 1'b0;
    wire _936 = 1'b0;
    wire _935 = 1'b0;
    wire _933 = 1'b0;
    wire _932 = 1'b0;
    wire _930 = 1'b0;
    wire _929 = 1'b0;
    wire _927 = 1'b0;
    wire _926 = 1'b0;
    wire _924 = 1'b0;
    wire _923 = 1'b0;
    wire _921 = 1'b0;
    wire _920 = 1'b0;
    wire _918 = 1'b0;
    wire _917 = 1'b0;
    reg _919;
    reg _922;
    reg _925;
    reg _928;
    reg _931;
    reg _934;
    reg _937;
    reg _940;
    reg _943;
    wire _944;
    wire _915 = 1'b0;
    wire _914 = 1'b0;
    wire _912 = 1'b0;
    wire _911 = 1'b0;
    wire _909 = 1'b0;
    wire _908 = 1'b0;
    wire _906 = 1'b0;
    wire _905 = 1'b0;
    wire _903 = 1'b0;
    wire _902 = 1'b0;
    wire _900 = 1'b0;
    wire _899 = 1'b0;
    wire _897 = 1'b0;
    wire _896 = 1'b0;
    wire _894 = 1'b0;
    wire _893 = 1'b0;
    wire _891 = 1'b0;
    wire _890 = 1'b0;
    reg _892;
    reg _895;
    reg _898;
    reg _901;
    reg _904;
    reg _907;
    reg _910;
    reg _913;
    reg _916;
    wire _945;
    wire _946;
    wire write_enable_46;
    wire _951;
    wire [131:0] _958;
    wire [63:0] _959;
    wire _887 = 1'b0;
    wire _886 = 1'b0;
    wire _889;
    wire _31;
    reg PHASE_10;
    wire [63:0] _971;
    wire [11:0] address_47;
    wire write_enable_47;
    wire [11:0] address_48;
    wire _1158;
    wire read_enable_39;
    wire _1156;
    wire write_enable_48;
    wire _1160;
    wire [131:0] _1165;
    wire [63:0] _1166;
    wire [11:0] _1151 = 12'b000000000000;
    wire [11:0] address_49;
    wire _1149;
    wire write_enable_49;
    wire [63:0] _1074;
    wire [63:0] _1073;
    wire [63:0] _1075;
    wire [63:0] _1071;
    wire [63:0] _1070;
    wire [63:0] q1_3;
    wire [63:0] _1076;
    wire [11:0] address_50;
    wire write_enable_50 = 1'b0;
    wire _1061;
    wire read_enable_40;
    wire [11:0] address_51;
    wire _1057;
    wire read_enable_41;
    wire _1055;
    wire write_enable_51;
    wire _1059;
    wire [131:0] _1066;
    wire [63:0] _1067;
    wire [63:0] data_47 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_48;
    wire [11:0] _1049 = 12'b000000000000;
    wire _1047;
    wire _1046;
    wire _1045;
    wire _1044;
    wire _1043;
    wire _1042;
    wire _1041;
    wire _1040;
    wire _1039;
    wire _1038;
    wire _1037;
    wire _1036;
    wire [11:0] _1048;
    wire [11:0] address_52;
    wire write_enable_52 = 1'b0;
    wire _1033;
    wire read_enable_42;
    wire [63:0] data_49;
    wire [63:0] data_50;
    wire _1030;
    wire _1029;
    wire _1028;
    wire _1027;
    wire _1026;
    wire _1025;
    wire _1024;
    wire _1023;
    wire _1022;
    wire _1021;
    wire _1020;
    wire _1019;
    wire [11:0] _1031;
    wire [11:0] address_53;
    wire _1016;
    wire read_enable_43;
    wire _1014;
    wire write_enable_53;
    wire _1018;
    wire [131:0] _1053;
    wire [63:0] _1054;
    wire _973 = 1'b0;
    wire _972 = 1'b0;
    wire _975;
    wire _35;
    reg PHASE_11;
    wire [63:0] _1068;
    wire [11:0] address_54;
    wire _1006;
    wire read_enable_44;
    wire write_enable_54;
    wire _1008;
    wire [11:0] address_55;
    wire _1001;
    wire read_enable_45;
    wire _999;
    wire write_enable_55;
    wire _1003;
    wire [131:0] _1011;
    wire [63:0] _1012;
    wire [63:0] _1079;
    wire [63:0] data_51;
    wire [63:0] data_52;
    wire [63:0] data_53;
    wire [63:0] data_54;
    wire [11:0] address_56;
    wire _992;
    wire read_enable_46;
    wire _989;
    wire _990;
    wire write_enable_56;
    wire _994;
    wire [11:0] address_57;
    wire _985;
    wire read_enable_47;
    wire _982;
    wire _983;
    wire write_enable_57;
    wire _987;
    wire [131:0] _997;
    wire [63:0] _998;
    wire _980 = 1'b0;
    wire _979 = 1'b0;
    wire _1080;
    wire _37;
    reg PHASE_12;
    wire [63:0] q0_3;
    wire _977 = 1'b0;
    wire _976 = 1'b0;
    reg _978;
    wire [63:0] _1069;
    wire [191:0] _1078;
    wire [63:0] _1081;
    wire [63:0] data_55;
    wire [63:0] data_56;
    wire [63:0] data_57;
    wire [63:0] data_58;
    wire [11:0] address_58;
    wire _1145;
    wire _1144;
    wire read_enable_48;
    wire _1138 = 1'b0;
    wire _1137 = 1'b0;
    wire _1135 = 1'b0;
    wire _1134 = 1'b0;
    wire _1132 = 1'b0;
    wire _1131 = 1'b0;
    wire _1129 = 1'b0;
    wire _1128 = 1'b0;
    wire _1126 = 1'b0;
    wire _1125 = 1'b0;
    wire _1123 = 1'b0;
    wire _1122 = 1'b0;
    wire _1120 = 1'b0;
    wire _1119 = 1'b0;
    wire _1117 = 1'b0;
    wire _1116 = 1'b0;
    wire _1114 = 1'b0;
    wire _1113 = 1'b0;
    reg _1115;
    reg _1118;
    reg _1121;
    reg _1124;
    reg _1127;
    reg _1130;
    reg _1133;
    reg _1136;
    reg _1139;
    wire _1140;
    wire _1111 = 1'b0;
    wire _1110 = 1'b0;
    wire _1108 = 1'b0;
    wire _1107 = 1'b0;
    wire _1105 = 1'b0;
    wire _1104 = 1'b0;
    wire _1102 = 1'b0;
    wire _1101 = 1'b0;
    wire _1099 = 1'b0;
    wire _1098 = 1'b0;
    wire _1096 = 1'b0;
    wire _1095 = 1'b0;
    wire _1093 = 1'b0;
    wire _1092 = 1'b0;
    wire _1090 = 1'b0;
    wire _1089 = 1'b0;
    wire _1087 = 1'b0;
    wire _1086 = 1'b0;
    reg _1088;
    reg _1091;
    reg _1094;
    reg _1097;
    reg _1100;
    reg _1103;
    reg _1106;
    reg _1109;
    reg _1112;
    wire _1141;
    wire _1142;
    wire write_enable_58;
    wire _1147;
    wire [131:0] _1154;
    wire [63:0] _1155;
    wire _1083 = 1'b0;
    wire _1082 = 1'b0;
    wire _1085;
    wire _39;
    reg PHASE_13;
    wire [63:0] _1167;
    wire [11:0] address_59;
    wire write_enable_59;
    wire [11:0] address_60;
    wire _1354;
    wire read_enable_49;
    wire _1352;
    wire write_enable_60;
    wire _1356;
    wire [131:0] _1361;
    wire [63:0] _1362;
    wire [11:0] _1347 = 12'b000000000000;
    wire [11:0] address_61;
    wire _1345;
    wire write_enable_61;
    wire [63:0] _1270;
    wire [63:0] _1269;
    wire [63:0] _1271;
    wire [63:0] _1267;
    wire [63:0] _1266;
    wire [63:0] q1_4;
    wire [63:0] _1272;
    wire [11:0] address_62;
    wire write_enable_62 = 1'b0;
    wire _1257;
    wire read_enable_50;
    wire [11:0] address_63;
    wire _1253;
    wire read_enable_51;
    wire _1251;
    wire write_enable_63;
    wire _1255;
    wire [131:0] _1262;
    wire [63:0] _1263;
    wire [63:0] data_59 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_60;
    wire [11:0] _1245 = 12'b000000000000;
    wire _1243;
    wire _1242;
    wire _1241;
    wire _1240;
    wire _1239;
    wire _1238;
    wire _1237;
    wire _1236;
    wire _1235;
    wire _1234;
    wire _1233;
    wire _1232;
    wire [11:0] _1244;
    wire [11:0] address_64;
    wire write_enable_64 = 1'b0;
    wire _1229;
    wire read_enable_52;
    wire [63:0] data_61;
    wire [63:0] data_62;
    wire _1226;
    wire _1225;
    wire _1224;
    wire _1223;
    wire _1222;
    wire _1221;
    wire _1220;
    wire _1219;
    wire _1218;
    wire _1217;
    wire _1216;
    wire _1215;
    wire [11:0] _1227;
    wire [11:0] address_65;
    wire _1212;
    wire read_enable_53;
    wire _1210;
    wire write_enable_65;
    wire _1214;
    wire [131:0] _1249;
    wire [63:0] _1250;
    wire _1169 = 1'b0;
    wire _1168 = 1'b0;
    wire _1171;
    wire _43;
    reg PHASE_14;
    wire [63:0] _1264;
    wire [11:0] address_66;
    wire _1202;
    wire read_enable_54;
    wire write_enable_66;
    wire _1204;
    wire [11:0] address_67;
    wire _1197;
    wire read_enable_55;
    wire _1195;
    wire write_enable_67;
    wire _1199;
    wire [131:0] _1207;
    wire [63:0] _1208;
    wire [63:0] _1275;
    wire [63:0] data_63;
    wire [63:0] data_64;
    wire [63:0] data_65;
    wire [63:0] data_66;
    wire [11:0] address_68;
    wire _1188;
    wire read_enable_56;
    wire _1185;
    wire _1186;
    wire write_enable_68;
    wire _1190;
    wire [11:0] address_69;
    wire _1181;
    wire read_enable_57;
    wire _1178;
    wire _1179;
    wire write_enable_69;
    wire _1183;
    wire [131:0] _1193;
    wire [63:0] _1194;
    wire _1176 = 1'b0;
    wire _1175 = 1'b0;
    wire _1276;
    wire _45;
    reg PHASE_15;
    wire [63:0] q0_4;
    wire _1173 = 1'b0;
    wire _1172 = 1'b0;
    reg _1174;
    wire [63:0] _1265;
    wire [191:0] _1274;
    wire [63:0] _1277;
    wire [63:0] data_67;
    wire [63:0] data_68;
    wire [63:0] data_69;
    wire [63:0] data_70;
    wire [11:0] address_70;
    wire _1341;
    wire _1340;
    wire read_enable_58;
    wire _1334 = 1'b0;
    wire _1333 = 1'b0;
    wire _1331 = 1'b0;
    wire _1330 = 1'b0;
    wire _1328 = 1'b0;
    wire _1327 = 1'b0;
    wire _1325 = 1'b0;
    wire _1324 = 1'b0;
    wire _1322 = 1'b0;
    wire _1321 = 1'b0;
    wire _1319 = 1'b0;
    wire _1318 = 1'b0;
    wire _1316 = 1'b0;
    wire _1315 = 1'b0;
    wire _1313 = 1'b0;
    wire _1312 = 1'b0;
    wire _1310 = 1'b0;
    wire _1309 = 1'b0;
    reg _1311;
    reg _1314;
    reg _1317;
    reg _1320;
    reg _1323;
    reg _1326;
    reg _1329;
    reg _1332;
    reg _1335;
    wire _1336;
    wire _1307 = 1'b0;
    wire _1306 = 1'b0;
    wire _1304 = 1'b0;
    wire _1303 = 1'b0;
    wire _1301 = 1'b0;
    wire _1300 = 1'b0;
    wire _1298 = 1'b0;
    wire _1297 = 1'b0;
    wire _1295 = 1'b0;
    wire _1294 = 1'b0;
    wire _1292 = 1'b0;
    wire _1291 = 1'b0;
    wire _1289 = 1'b0;
    wire _1288 = 1'b0;
    wire _1286 = 1'b0;
    wire _1285 = 1'b0;
    wire _1283 = 1'b0;
    wire _1282 = 1'b0;
    reg _1284;
    reg _1287;
    reg _1290;
    reg _1293;
    reg _1296;
    reg _1299;
    reg _1302;
    reg _1305;
    reg _1308;
    wire _1337;
    wire _1338;
    wire write_enable_70;
    wire _1343;
    wire [131:0] _1350;
    wire [63:0] _1351;
    wire _1279 = 1'b0;
    wire _1278 = 1'b0;
    wire _1281;
    wire _47;
    reg PHASE_16;
    wire [63:0] _1363;
    wire [11:0] address_71;
    wire write_enable_71;
    wire [11:0] address_72;
    wire _1550;
    wire read_enable_59;
    wire _1548;
    wire write_enable_72;
    wire _1552;
    wire [131:0] _1557;
    wire [63:0] _1558;
    wire [11:0] _1543 = 12'b000000000000;
    wire [11:0] address_73;
    wire _1541;
    wire write_enable_73;
    wire [63:0] _1466;
    wire [63:0] _1465;
    wire [63:0] _1467;
    wire [63:0] _1463;
    wire [63:0] _1462;
    wire [63:0] q1_5;
    wire [63:0] _1468;
    wire [11:0] address_74;
    wire write_enable_74 = 1'b0;
    wire _1453;
    wire read_enable_60;
    wire [11:0] address_75;
    wire _1449;
    wire read_enable_61;
    wire _1447;
    wire write_enable_75;
    wire _1451;
    wire [131:0] _1458;
    wire [63:0] _1459;
    wire [63:0] data_71 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_72;
    wire [11:0] _1441 = 12'b000000000000;
    wire _1439;
    wire _1438;
    wire _1437;
    wire _1436;
    wire _1435;
    wire _1434;
    wire _1433;
    wire _1432;
    wire _1431;
    wire _1430;
    wire _1429;
    wire _1428;
    wire [11:0] _1440;
    wire [11:0] address_76;
    wire write_enable_76 = 1'b0;
    wire _1425;
    wire read_enable_62;
    wire [63:0] data_73;
    wire [63:0] data_74;
    wire _1422;
    wire _1421;
    wire _1420;
    wire _1419;
    wire _1418;
    wire _1417;
    wire _1416;
    wire _1415;
    wire _1414;
    wire _1413;
    wire _1412;
    wire _1411;
    wire [11:0] _1423;
    wire [11:0] address_77;
    wire _1408;
    wire read_enable_63;
    wire _1406;
    wire write_enable_77;
    wire _1410;
    wire [131:0] _1445;
    wire [63:0] _1446;
    wire _1365 = 1'b0;
    wire _1364 = 1'b0;
    wire _1367;
    wire _51;
    reg PHASE_17;
    wire [63:0] _1460;
    wire [11:0] address_78;
    wire _1398;
    wire read_enable_64;
    wire write_enable_78;
    wire _1400;
    wire [11:0] address_79;
    wire _1393;
    wire read_enable_65;
    wire _1391;
    wire write_enable_79;
    wire _1395;
    wire [131:0] _1403;
    wire [63:0] _1404;
    wire [63:0] _1471;
    wire [63:0] data_75;
    wire [63:0] data_76;
    wire [63:0] data_77;
    wire [63:0] data_78;
    wire [11:0] address_80;
    wire _1384;
    wire read_enable_66;
    wire _1381;
    wire _1382;
    wire write_enable_80;
    wire _1386;
    wire [11:0] address_81;
    wire _1377;
    wire read_enable_67;
    wire _1374;
    wire _1375;
    wire write_enable_81;
    wire _1379;
    wire [131:0] _1389;
    wire [63:0] _1390;
    wire _1372 = 1'b0;
    wire _1371 = 1'b0;
    wire _1472;
    wire _53;
    reg PHASE_18;
    wire [63:0] q0_5;
    wire _1369 = 1'b0;
    wire _1368 = 1'b0;
    reg _1370;
    wire [63:0] _1461;
    wire [191:0] _1470;
    wire [63:0] _1473;
    wire [63:0] data_79;
    wire [63:0] data_80;
    wire [63:0] data_81;
    wire [63:0] data_82;
    wire [11:0] address_82;
    wire _1537;
    wire _1536;
    wire read_enable_68;
    wire _1530 = 1'b0;
    wire _1529 = 1'b0;
    wire _1527 = 1'b0;
    wire _1526 = 1'b0;
    wire _1524 = 1'b0;
    wire _1523 = 1'b0;
    wire _1521 = 1'b0;
    wire _1520 = 1'b0;
    wire _1518 = 1'b0;
    wire _1517 = 1'b0;
    wire _1515 = 1'b0;
    wire _1514 = 1'b0;
    wire _1512 = 1'b0;
    wire _1511 = 1'b0;
    wire _1509 = 1'b0;
    wire _1508 = 1'b0;
    wire _1506 = 1'b0;
    wire _1505 = 1'b0;
    reg _1507;
    reg _1510;
    reg _1513;
    reg _1516;
    reg _1519;
    reg _1522;
    reg _1525;
    reg _1528;
    reg _1531;
    wire _1532;
    wire _1503 = 1'b0;
    wire _1502 = 1'b0;
    wire _1500 = 1'b0;
    wire _1499 = 1'b0;
    wire _1497 = 1'b0;
    wire _1496 = 1'b0;
    wire _1494 = 1'b0;
    wire _1493 = 1'b0;
    wire _1491 = 1'b0;
    wire _1490 = 1'b0;
    wire _1488 = 1'b0;
    wire _1487 = 1'b0;
    wire _1485 = 1'b0;
    wire _1484 = 1'b0;
    wire _1482 = 1'b0;
    wire _1481 = 1'b0;
    wire _1479 = 1'b0;
    wire _1478 = 1'b0;
    reg _1480;
    reg _1483;
    reg _1486;
    reg _1489;
    reg _1492;
    reg _1495;
    reg _1498;
    reg _1501;
    reg _1504;
    wire _1533;
    wire _1534;
    wire write_enable_82;
    wire _1539;
    wire [131:0] _1546;
    wire [63:0] _1547;
    wire _1475 = 1'b0;
    wire _1474 = 1'b0;
    wire _1477;
    wire _55;
    reg PHASE_19;
    wire [63:0] _1559;
    wire [11:0] address_83;
    wire write_enable_83;
    wire [11:0] address_84;
    wire _1746;
    wire read_enable_69;
    wire _1744;
    wire write_enable_84;
    wire _1748;
    wire [131:0] _1753;
    wire [63:0] _1754;
    wire [11:0] _1739 = 12'b000000000000;
    wire [11:0] address_85;
    wire _1737;
    wire write_enable_85;
    wire [3:0] _292;
    wire _291;
    wire _289;
    wire [63:0] _288;
    wire [63:0] _287;
    wire [63:0] _286;
    wire [63:0] _285;
    wire [63:0] _284;
    wire [63:0] _283;
    wire [63:0] _282;
    wire [63:0] _1662;
    wire [63:0] _1661;
    wire [63:0] _1663;
    wire [63:0] _1659;
    wire [63:0] _1658;
    wire [63:0] q1_6;
    wire [63:0] _1664;
    wire [11:0] address_86;
    wire write_enable_86 = 1'b0;
    wire _1649;
    wire read_enable_70;
    wire [11:0] address_87;
    wire _1645;
    wire read_enable_71;
    wire _1643;
    wire write_enable_87;
    wire _1647;
    wire [131:0] _1654;
    wire [63:0] _1655;
    wire [63:0] data_83 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] data_84;
    wire [11:0] _1637 = 12'b000000000000;
    wire _1635;
    wire _1634;
    wire _1633;
    wire _1632;
    wire _1631;
    wire _1630;
    wire _1629;
    wire _1628;
    wire _1627;
    wire _1626;
    wire _1625;
    wire _1624;
    wire [11:0] _1636;
    wire [11:0] address_88;
    wire write_enable_88 = 1'b0;
    wire _1621;
    wire read_enable_72;
    wire [63:0] data_85;
    wire [63:0] data_86;
    wire [11:0] _60;
    wire _1618;
    wire _1617;
    wire _1616;
    wire _1615;
    wire _1614;
    wire _1613;
    wire _1612;
    wire _1611;
    wire _1610;
    wire _1609;
    wire _1608;
    wire _1607;
    wire [11:0] _1619;
    wire [11:0] address_89;
    wire _1604;
    wire read_enable_73;
    wire [7:0] _62;
    wire _1602;
    wire write_enable_89;
    wire _1606;
    wire [131:0] _1641;
    wire [63:0] _1642;
    wire _1561 = 1'b0;
    wire _1560 = 1'b0;
    wire _1563;
    wire _63;
    reg PHASE_20;
    wire [63:0] _1656;
    wire [11:0] address_90;
    wire _1594;
    wire read_enable_74;
    wire write_enable_90;
    wire _1596;
    wire [11:0] address_91;
    wire _1589;
    wire read_enable_75;
    wire _1587;
    wire write_enable_91;
    wire _1591;
    wire [131:0] _1599;
    wire [63:0] _1600;
    wire [63:0] _1667;
    wire [63:0] data_87;
    wire [63:0] data_88;
    wire [63:0] data_89;
    wire [63:0] data_90;
    wire [11:0] _198 = 12'b000000000000;
    wire [11:0] _197 = 12'b000000000000;
    wire [11:0] _195 = 12'b000000000000;
    wire [11:0] _194 = 12'b000000000000;
    wire [11:0] _192 = 12'b000000000000;
    wire [11:0] _191 = 12'b000000000000;
    wire [11:0] _189 = 12'b000000000000;
    wire [11:0] _188 = 12'b000000000000;
    wire [11:0] _186 = 12'b000000000000;
    wire [11:0] _185 = 12'b000000000000;
    wire [11:0] _183 = 12'b000000000000;
    wire [11:0] _182 = 12'b000000000000;
    wire [11:0] _180 = 12'b000000000000;
    wire [11:0] _179 = 12'b000000000000;
    wire [11:0] _177 = 12'b000000000000;
    wire [11:0] _176 = 12'b000000000000;
    wire [11:0] _174 = 12'b000000000000;
    wire [11:0] _173 = 12'b000000000000;
    reg [11:0] _175;
    reg [11:0] _178;
    reg [11:0] _181;
    reg [11:0] _184;
    reg [11:0] _187;
    reg [11:0] _190;
    reg [11:0] _193;
    reg [11:0] _196;
    reg [11:0] _199;
    wire [11:0] _172;
    wire [11:0] address_92;
    wire _1580;
    wire read_enable_76;
    wire _1577;
    wire _1578;
    wire write_enable_92;
    wire _1582;
    wire [11:0] address_93;
    wire _1573;
    wire read_enable_77;
    wire _1570;
    wire _1571;
    wire write_enable_93;
    wire _1575;
    wire [131:0] _1585;
    wire [63:0] _1586;
    wire _99;
    wire _1568 = 1'b0;
    wire _1567 = 1'b0;
    wire _1668;
    wire _65;
    reg PHASE_21;
    wire [63:0] q0_6;
    wire _1565 = 1'b0;
    wire _1564 = 1'b0;
    wire _92;
    reg _1566;
    wire [63:0] _1657;
    wire [191:0] _1666;
    wire [63:0] _1669;
    wire [63:0] data_91;
    wire [63:0] data_92;
    wire [63:0] data_93;
    wire [63:0] data_94;
    wire [11:0] _163 = 12'b000000000000;
    wire [11:0] _162 = 12'b000000000000;
    wire [11:0] _160 = 12'b000000000000;
    wire [11:0] _159 = 12'b000000000000;
    wire [11:0] _157 = 12'b000000000000;
    wire [11:0] _156 = 12'b000000000000;
    wire [11:0] _154 = 12'b000000000000;
    wire [11:0] _153 = 12'b000000000000;
    wire [11:0] _151 = 12'b000000000000;
    wire [11:0] _150 = 12'b000000000000;
    wire [11:0] _148 = 12'b000000000000;
    wire [11:0] _147 = 12'b000000000000;
    wire [11:0] _145 = 12'b000000000000;
    wire [11:0] _144 = 12'b000000000000;
    wire [11:0] _142 = 12'b000000000000;
    wire [11:0] _141 = 12'b000000000000;
    wire [11:0] _139 = 12'b000000000000;
    wire [11:0] _138 = 12'b000000000000;
    wire [11:0] _137;
    reg [11:0] _140;
    reg [11:0] _143;
    reg [11:0] _146;
    reg [11:0] _149;
    reg [11:0] _152;
    reg [11:0] _155;
    reg [11:0] _158;
    reg [11:0] _161;
    reg [11:0] _164;
    wire [11:0] _68;
    wire [11:0] address_94;
    wire _1733;
    wire [7:0] _70;
    wire _1732;
    wire read_enable_78;
    wire _1726 = 1'b0;
    wire _1725 = 1'b0;
    wire _1723 = 1'b0;
    wire _1722 = 1'b0;
    wire _1720 = 1'b0;
    wire _1719 = 1'b0;
    wire _1717 = 1'b0;
    wire _1716 = 1'b0;
    wire _1714 = 1'b0;
    wire _1713 = 1'b0;
    wire _1711 = 1'b0;
    wire _1710 = 1'b0;
    wire _1708 = 1'b0;
    wire _1707 = 1'b0;
    wire _1705 = 1'b0;
    wire _1704 = 1'b0;
    wire _1702 = 1'b0;
    wire _1701 = 1'b0;
    wire _290;
    reg _1703;
    reg _1706;
    reg _1709;
    reg _1712;
    reg _1715;
    reg _1718;
    reg _1721;
    reg _1724;
    reg _1727;
    wire _1728;
    wire _1699 = 1'b0;
    wire _1698 = 1'b0;
    wire _1696 = 1'b0;
    wire _1695 = 1'b0;
    wire _1693 = 1'b0;
    wire _1692 = 1'b0;
    wire _1690 = 1'b0;
    wire _1689 = 1'b0;
    wire _1687 = 1'b0;
    wire _1686 = 1'b0;
    wire _1684 = 1'b0;
    wire _1683 = 1'b0;
    wire _1681 = 1'b0;
    wire _1680 = 1'b0;
    wire _1678 = 1'b0;
    wire _1677 = 1'b0;
    wire _1675 = 1'b0;
    wire _1674 = 1'b0;
    wire _130;
    reg _1676;
    reg _1679;
    reg _1682;
    reg _1685;
    reg _1688;
    reg _1691;
    reg _1694;
    reg _1697;
    reg _1700;
    wire _1729;
    wire _128 = 1'b0;
    wire _127 = 1'b0;
    wire _125 = 1'b0;
    wire _124 = 1'b0;
    wire _122 = 1'b0;
    wire _121 = 1'b0;
    wire _119 = 1'b0;
    wire _118 = 1'b0;
    wire _116 = 1'b0;
    wire _115 = 1'b0;
    wire _113 = 1'b0;
    wire _112 = 1'b0;
    wire _110 = 1'b0;
    wire _109 = 1'b0;
    wire _107 = 1'b0;
    wire _106 = 1'b0;
    wire vdd = 1'b1;
    wire _104 = 1'b0;
    wire _103 = 1'b0;
    wire _102;
    reg _105;
    reg _108;
    reg _111;
    reg _114;
    reg _117;
    reg _120;
    reg _123;
    reg _126;
    reg _129;
    wire _1730;
    wire write_enable_94;
    wire _1735;
    wire gnd = 1'b0;
    wire [131:0] _1742;
    wire [63:0] _1743;
    wire _72;
    wire _1671 = 1'b0;
    wire _1670 = 1'b0;
    wire _1673;
    wire _73;
    reg PHASE_22;
    wire [63:0] _1755;
    wire _76;
    wire _78;
    wire _80;
    wire _82;
    wire _84;
    wire [523:0] _91;
    wire _1756;

    /* logic */
    assign address = _372 ? _199 : _367;
    assign write_enable = _365 & _372;
    assign address_0 = _372 ? _164 : _68;
    assign _374 = ~ _372;
    assign read_enable = _360 & _374;
    assign _372 = ~ PHASE_1;
    assign write_enable_0 = _358 & _372;
    assign _376 = write_enable_0 | read_enable;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_376), .regcea(vdd), .wea(write_enable_0), .addra(address_0), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable), .regceb(vdd), .web(write_enable), .addrb(address), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_381[131:131]), .sbiterrb(_381[130:130]), .doutb(_381[129:66]), .dbiterra(_381[65:65]), .sbiterra(_381[64:64]), .douta(_381[63:0]) );
    assign _382 = _381[63:0];
    assign address_1 = PHASE_1 ? _199 : _367;
    assign _365 = _129 & _328;
    assign write_enable_1 = _365 & PHASE_1;
    assign _279 = _271[129:66];
    assign _278 = _258[129:66];
    assign _280 = PHASE ? _279 : _278;
    assign _276 = _216[129:66];
    assign _275 = _202[129:66];
    assign q1 = PHASE_0 ? _276 : _275;
    assign _281 = _96 ? _280 : q1;
    assign address_2 = _260 ? _254 : _253;
    assign _266 = ~ _260;
    assign read_enable_0 = _102 & _266;
    assign address_3 = _260 ? _60 : _236;
    assign _262 = ~ _260;
    assign read_enable_1 = _102 & _262;
    assign _260 = ~ PHASE;
    assign write_enable_3 = _219 & _260;
    assign _264 = write_enable_3 | read_enable_1;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_0
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_264), .regcea(vdd), .wea(write_enable_3), .addra(address_3), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_0), .regceb(vdd), .web(write_enable_2), .addrb(address_2), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_271[131:131]), .sbiterrb(_271[130:130]), .doutb(_271[129:66]), .dbiterra(_271[65:65]), .sbiterra(_271[64:64]), .douta(_271[63:0]) );
    assign _272 = _271[63:0];
    assign _252 = _172[11:11];
    assign _251 = _172[10:10];
    assign _250 = _172[9:9];
    assign _249 = _172[8:8];
    assign _248 = _172[7:7];
    assign _247 = _172[6:6];
    assign _246 = _172[5:5];
    assign _245 = _172[4:4];
    assign _244 = _172[3:3];
    assign _243 = _172[2:2];
    assign _242 = _172[1:1];
    assign _241 = _172[0:0];
    assign _253 = { _241, _242, _243, _244, _245, _246, _247, _248, _249, _250, _251, _252 };
    assign address_4 = PHASE ? _254 : _253;
    assign _238 = ~ PHASE;
    assign read_enable_2 = _102 & _238;
    assign data_1 = wr_d7;
    assign _235 = _137[11:11];
    assign _234 = _137[10:10];
    assign _233 = _137[9:9];
    assign _232 = _137[8:8];
    assign _231 = _137[7:7];
    assign _230 = _137[6:6];
    assign _229 = _137[5:5];
    assign _228 = _137[4:4];
    assign _227 = _137[3:3];
    assign _226 = _137[2:2];
    assign _225 = _137[1:1];
    assign _224 = _137[0:0];
    assign _236 = { _224, _225, _226, _227, _228, _229, _230, _231, _232, _233, _234, _235 };
    assign address_5 = PHASE ? _60 : _236;
    assign _221 = ~ PHASE;
    assign read_enable_3 = _102 & _221;
    assign _219 = _62[7:7];
    assign write_enable_5 = _219 & PHASE;
    assign _223 = write_enable_5 | read_enable_3;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_1
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_223), .regcea(vdd), .wea(write_enable_5), .addra(address_5), .dina(data_1), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_2), .regceb(vdd), .web(write_enable_4), .addrb(address_4), .dinb(data), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_258[131:131]), .sbiterrb(_258[130:130]), .doutb(_258[129:66]), .dbiterra(_258[65:65]), .sbiterra(_258[64:64]), .douta(_258[63:0]) );
    assign _259 = _258[63:0];
    assign _89 = ~ PHASE;
    assign _3 = _89;
    always @(posedge _84) begin
        if (_82)
            PHASE <= _87;
        else
            if (_72)
                PHASE <= _3;
    end
    assign _273 = PHASE ? _272 : _259;
    assign address_6 = _204 ? _199 : _172;
    assign _211 = ~ _204;
    assign read_enable_4 = _102 & _211;
    assign write_enable_6 = _167 & _204;
    assign _213 = write_enable_6 | read_enable_4;
    assign address_7 = _204 ? _164 : _137;
    assign _206 = ~ _204;
    assign read_enable_5 = _102 & _206;
    assign _204 = ~ PHASE_0;
    assign write_enable_7 = _132 & _204;
    assign _208 = write_enable_7 | read_enable_5;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_2
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_208), .regcea(vdd), .wea(write_enable_7), .addra(address_7), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_213), .regceb(vdd), .web(write_enable_6), .addrb(address_6), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_216[131:131]), .sbiterrb(_216[130:130]), .doutb(_216[129:66]), .dbiterra(_216[65:65]), .sbiterra(_216[64:64]), .douta(_216[63:0]) );
    assign _217 = _216[63:0];
    assign _295 = _294[127:64];
    assign data_3 = _295;
    assign address_8 = PHASE_0 ? _199 : _172;
    assign _169 = ~ PHASE_0;
    assign read_enable_6 = _102 & _169;
    assign _166 = ~ _130;
    assign _167 = _129 & _166;
    assign write_enable_8 = _167 & PHASE_0;
    assign _171 = write_enable_8 | read_enable_6;
    assign address_9 = PHASE_0 ? _164 : _137;
    assign _134 = ~ PHASE_0;
    assign read_enable_7 = _102 & _134;
    assign _131 = ~ _130;
    assign _132 = _129 & _131;
    assign write_enable_9 = _132 & PHASE_0;
    assign _136 = write_enable_9 | read_enable_7;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_3
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_136), .regcea(vdd), .wea(write_enable_9), .addra(address_9), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_171), .regceb(vdd), .web(write_enable_8), .addrb(address_8), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_202[131:131]), .sbiterrb(_202[130:130]), .doutb(_202[129:66]), .dbiterra(_202[65:65]), .sbiterra(_202[64:64]), .douta(_202[63:0]) );
    assign _203 = _202[63:0];
    assign _296 = ~ PHASE_0;
    assign _5 = _296;
    always @(posedge _84) begin
        if (_82)
            PHASE_0 <= _98;
        else
            if (_99)
                PHASE_0 <= _5;
    end
    assign q0 = PHASE_0 ? _217 : _203;
    always @(posedge _84) begin
        if (_82)
            _96 <= _94;
        else
            _96 <= _92;
    end
    assign _274 = _96 ? _273 : q0;
    dp_62
        dp_6
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_274), .d2(_281), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_294[191:128]), .q2(_294[127:64]), .q1(_294[63:0]) );
    assign _297 = _294[63:0];
    assign data_7 = _297;
    assign address_10 = PHASE_1 ? _164 : _68;
    assign _361 = ~ PHASE_1;
    assign _360 = _70[7:7];
    assign read_enable_8 = _360 & _361;
    always @(posedge _84) begin
        if (_82)
            _331 <= _330;
        else
            _331 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _334 <= _333;
        else
            _334 <= _331;
    end
    always @(posedge _84) begin
        if (_82)
            _337 <= _336;
        else
            _337 <= _334;
    end
    always @(posedge _84) begin
        if (_82)
            _340 <= _339;
        else
            _340 <= _337;
    end
    always @(posedge _84) begin
        if (_82)
            _343 <= _342;
        else
            _343 <= _340;
    end
    always @(posedge _84) begin
        if (_82)
            _346 <= _345;
        else
            _346 <= _343;
    end
    always @(posedge _84) begin
        if (_82)
            _349 <= _348;
        else
            _349 <= _346;
    end
    always @(posedge _84) begin
        if (_82)
            _352 <= _351;
        else
            _352 <= _349;
    end
    always @(posedge _84) begin
        if (_82)
            _355 <= _354;
        else
            _355 <= _352;
    end
    assign _356 = ~ _355;
    always @(posedge _84) begin
        if (_82)
            _304 <= _303;
        else
            _304 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _307 <= _306;
        else
            _307 <= _304;
    end
    always @(posedge _84) begin
        if (_82)
            _310 <= _309;
        else
            _310 <= _307;
    end
    always @(posedge _84) begin
        if (_82)
            _313 <= _312;
        else
            _313 <= _310;
    end
    always @(posedge _84) begin
        if (_82)
            _316 <= _315;
        else
            _316 <= _313;
    end
    always @(posedge _84) begin
        if (_82)
            _319 <= _318;
        else
            _319 <= _316;
    end
    always @(posedge _84) begin
        if (_82)
            _322 <= _321;
        else
            _322 <= _319;
    end
    always @(posedge _84) begin
        if (_82)
            _325 <= _324;
        else
            _325 <= _322;
    end
    always @(posedge _84) begin
        if (_82)
            _328 <= _327;
        else
            _328 <= _325;
    end
    assign _357 = _328 & _356;
    assign _358 = _129 & _357;
    assign write_enable_10 = _358 & PHASE_1;
    assign _363 = write_enable_10 | read_enable_8;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_4
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_363), .regcea(vdd), .wea(write_enable_10), .addra(address_10), .dina(data_7), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_1), .regceb(vdd), .web(write_enable_1), .addrb(address_1), .dinb(data_3), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_370[131:131]), .sbiterrb(_370[130:130]), .doutb(_370[129:66]), .dbiterra(_370[65:65]), .sbiterra(_370[64:64]), .douta(_370[63:0]) );
    assign _371 = _370[63:0];
    assign _301 = ~ PHASE_1;
    assign _7 = _301;
    always @(posedge _84) begin
        if (_82)
            PHASE_1 <= _299;
        else
            if (_72)
                PHASE_1 <= _7;
    end
    assign _383 = PHASE_1 ? _382 : _371;
    assign address_11 = _568 ? _199 : _563;
    assign write_enable_11 = _561 & _568;
    assign address_12 = _568 ? _164 : _68;
    assign _570 = ~ _568;
    assign read_enable_9 = _556 & _570;
    assign _568 = ~ PHASE_4;
    assign write_enable_12 = _554 & _568;
    assign _572 = write_enable_12 | read_enable_9;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_5
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_572), .regcea(vdd), .wea(write_enable_12), .addra(address_12), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_11), .regceb(vdd), .web(write_enable_11), .addrb(address_11), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_577[131:131]), .sbiterrb(_577[130:130]), .doutb(_577[129:66]), .dbiterra(_577[65:65]), .sbiterra(_577[64:64]), .douta(_577[63:0]) );
    assign _578 = _577[63:0];
    assign address_13 = PHASE_4 ? _199 : _563;
    assign _561 = _129 & _524;
    assign write_enable_13 = _561 & PHASE_4;
    assign _486 = _478[129:66];
    assign _485 = _465[129:66];
    assign _487 = PHASE_2 ? _486 : _485;
    assign _483 = _423[129:66];
    assign _482 = _409[129:66];
    assign q1_0 = PHASE_3 ? _483 : _482;
    assign _488 = _390 ? _487 : q1_0;
    assign address_14 = _467 ? _461 : _460;
    assign _473 = ~ _467;
    assign read_enable_10 = _102 & _473;
    assign address_15 = _467 ? _60 : _443;
    assign _469 = ~ _467;
    assign read_enable_11 = _102 & _469;
    assign _467 = ~ PHASE_2;
    assign write_enable_15 = _426 & _467;
    assign _471 = write_enable_15 | read_enable_11;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_6
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_471), .regcea(vdd), .wea(write_enable_15), .addra(address_15), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_10), .regceb(vdd), .web(write_enable_14), .addrb(address_14), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_478[131:131]), .sbiterrb(_478[130:130]), .doutb(_478[129:66]), .dbiterra(_478[65:65]), .sbiterra(_478[64:64]), .douta(_478[63:0]) );
    assign _479 = _478[63:0];
    assign _459 = _172[11:11];
    assign _458 = _172[10:10];
    assign _457 = _172[9:9];
    assign _456 = _172[8:8];
    assign _455 = _172[7:7];
    assign _454 = _172[6:6];
    assign _453 = _172[5:5];
    assign _452 = _172[4:4];
    assign _451 = _172[3:3];
    assign _450 = _172[2:2];
    assign _449 = _172[1:1];
    assign _448 = _172[0:0];
    assign _460 = { _448, _449, _450, _451, _452, _453, _454, _455, _456, _457, _458, _459 };
    assign address_16 = PHASE_2 ? _461 : _460;
    assign _445 = ~ PHASE_2;
    assign read_enable_12 = _102 & _445;
    assign data_13 = wr_d6;
    assign _442 = _137[11:11];
    assign _441 = _137[10:10];
    assign _440 = _137[9:9];
    assign _439 = _137[8:8];
    assign _438 = _137[7:7];
    assign _437 = _137[6:6];
    assign _436 = _137[5:5];
    assign _435 = _137[4:4];
    assign _434 = _137[3:3];
    assign _433 = _137[2:2];
    assign _432 = _137[1:1];
    assign _431 = _137[0:0];
    assign _443 = { _431, _432, _433, _434, _435, _436, _437, _438, _439, _440, _441, _442 };
    assign address_17 = PHASE_2 ? _60 : _443;
    assign _428 = ~ PHASE_2;
    assign read_enable_13 = _102 & _428;
    assign _426 = _62[6:6];
    assign write_enable_17 = _426 & PHASE_2;
    assign _430 = write_enable_17 | read_enable_13;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_7
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_430), .regcea(vdd), .wea(write_enable_17), .addra(address_17), .dina(data_13), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_12), .regceb(vdd), .web(write_enable_16), .addrb(address_16), .dinb(data_11), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_465[131:131]), .sbiterrb(_465[130:130]), .doutb(_465[129:66]), .dbiterra(_465[65:65]), .sbiterra(_465[64:64]), .douta(_465[63:0]) );
    assign _466 = _465[63:0];
    assign _387 = ~ PHASE_2;
    assign _11 = _387;
    always @(posedge _84) begin
        if (_82)
            PHASE_2 <= _385;
        else
            if (_72)
                PHASE_2 <= _11;
    end
    assign _480 = PHASE_2 ? _479 : _466;
    assign address_18 = _411 ? _199 : _172;
    assign _418 = ~ _411;
    assign read_enable_14 = _102 & _418;
    assign write_enable_18 = _402 & _411;
    assign _420 = write_enable_18 | read_enable_14;
    assign address_19 = _411 ? _164 : _137;
    assign _413 = ~ _411;
    assign read_enable_15 = _102 & _413;
    assign _411 = ~ PHASE_3;
    assign write_enable_19 = _395 & _411;
    assign _415 = write_enable_19 | read_enable_15;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_8
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_415), .regcea(vdd), .wea(write_enable_19), .addra(address_19), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_420), .regceb(vdd), .web(write_enable_18), .addrb(address_18), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_423[131:131]), .sbiterrb(_423[130:130]), .doutb(_423[129:66]), .dbiterra(_423[65:65]), .sbiterra(_423[64:64]), .douta(_423[63:0]) );
    assign _424 = _423[63:0];
    assign _491 = _490[127:64];
    assign data_15 = _491;
    assign address_20 = PHASE_3 ? _199 : _172;
    assign _404 = ~ PHASE_3;
    assign read_enable_16 = _102 & _404;
    assign _401 = ~ _130;
    assign _402 = _129 & _401;
    assign write_enable_20 = _402 & PHASE_3;
    assign _406 = write_enable_20 | read_enable_16;
    assign address_21 = PHASE_3 ? _164 : _137;
    assign _397 = ~ PHASE_3;
    assign read_enable_17 = _102 & _397;
    assign _394 = ~ _130;
    assign _395 = _129 & _394;
    assign write_enable_21 = _395 & PHASE_3;
    assign _399 = write_enable_21 | read_enable_17;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_9
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_399), .regcea(vdd), .wea(write_enable_21), .addra(address_21), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_406), .regceb(vdd), .web(write_enable_20), .addrb(address_20), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_409[131:131]), .sbiterrb(_409[130:130]), .doutb(_409[129:66]), .dbiterra(_409[65:65]), .sbiterra(_409[64:64]), .douta(_409[63:0]) );
    assign _410 = _409[63:0];
    assign _492 = ~ PHASE_3;
    assign _13 = _492;
    always @(posedge _84) begin
        if (_82)
            PHASE_3 <= _392;
        else
            if (_99)
                PHASE_3 <= _13;
    end
    assign q0_0 = PHASE_3 ? _424 : _410;
    always @(posedge _84) begin
        if (_82)
            _390 <= _389;
        else
            _390 <= _92;
    end
    assign _481 = _390 ? _480 : q0_0;
    dp_61
        dp_5
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_481), .d2(_488), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_490[191:128]), .q2(_490[127:64]), .q1(_490[63:0]) );
    assign _493 = _490[63:0];
    assign data_19 = _493;
    assign address_22 = PHASE_4 ? _164 : _68;
    assign _557 = ~ PHASE_4;
    assign _556 = _70[6:6];
    assign read_enable_18 = _556 & _557;
    always @(posedge _84) begin
        if (_82)
            _527 <= _526;
        else
            _527 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _530 <= _529;
        else
            _530 <= _527;
    end
    always @(posedge _84) begin
        if (_82)
            _533 <= _532;
        else
            _533 <= _530;
    end
    always @(posedge _84) begin
        if (_82)
            _536 <= _535;
        else
            _536 <= _533;
    end
    always @(posedge _84) begin
        if (_82)
            _539 <= _538;
        else
            _539 <= _536;
    end
    always @(posedge _84) begin
        if (_82)
            _542 <= _541;
        else
            _542 <= _539;
    end
    always @(posedge _84) begin
        if (_82)
            _545 <= _544;
        else
            _545 <= _542;
    end
    always @(posedge _84) begin
        if (_82)
            _548 <= _547;
        else
            _548 <= _545;
    end
    always @(posedge _84) begin
        if (_82)
            _551 <= _550;
        else
            _551 <= _548;
    end
    assign _552 = ~ _551;
    always @(posedge _84) begin
        if (_82)
            _500 <= _499;
        else
            _500 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _503 <= _502;
        else
            _503 <= _500;
    end
    always @(posedge _84) begin
        if (_82)
            _506 <= _505;
        else
            _506 <= _503;
    end
    always @(posedge _84) begin
        if (_82)
            _509 <= _508;
        else
            _509 <= _506;
    end
    always @(posedge _84) begin
        if (_82)
            _512 <= _511;
        else
            _512 <= _509;
    end
    always @(posedge _84) begin
        if (_82)
            _515 <= _514;
        else
            _515 <= _512;
    end
    always @(posedge _84) begin
        if (_82)
            _518 <= _517;
        else
            _518 <= _515;
    end
    always @(posedge _84) begin
        if (_82)
            _521 <= _520;
        else
            _521 <= _518;
    end
    always @(posedge _84) begin
        if (_82)
            _524 <= _523;
        else
            _524 <= _521;
    end
    assign _553 = _524 & _552;
    assign _554 = _129 & _553;
    assign write_enable_22 = _554 & PHASE_4;
    assign _559 = write_enable_22 | read_enable_18;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_10
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_559), .regcea(vdd), .wea(write_enable_22), .addra(address_22), .dina(data_19), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_13), .regceb(vdd), .web(write_enable_13), .addrb(address_13), .dinb(data_15), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_566[131:131]), .sbiterrb(_566[130:130]), .doutb(_566[129:66]), .dbiterra(_566[65:65]), .sbiterra(_566[64:64]), .douta(_566[63:0]) );
    assign _567 = _566[63:0];
    assign _497 = ~ PHASE_4;
    assign _15 = _497;
    always @(posedge _84) begin
        if (_82)
            PHASE_4 <= _495;
        else
            if (_72)
                PHASE_4 <= _15;
    end
    assign _579 = PHASE_4 ? _578 : _567;
    assign address_23 = _764 ? _199 : _759;
    assign write_enable_23 = _757 & _764;
    assign address_24 = _764 ? _164 : _68;
    assign _766 = ~ _764;
    assign read_enable_19 = _752 & _766;
    assign _764 = ~ PHASE_7;
    assign write_enable_24 = _750 & _764;
    assign _768 = write_enable_24 | read_enable_19;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_11
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_768), .regcea(vdd), .wea(write_enable_24), .addra(address_24), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_23), .regceb(vdd), .web(write_enable_23), .addrb(address_23), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_773[131:131]), .sbiterrb(_773[130:130]), .doutb(_773[129:66]), .dbiterra(_773[65:65]), .sbiterra(_773[64:64]), .douta(_773[63:0]) );
    assign _774 = _773[63:0];
    assign address_25 = PHASE_7 ? _199 : _759;
    assign _757 = _129 & _720;
    assign write_enable_25 = _757 & PHASE_7;
    assign _682 = _674[129:66];
    assign _681 = _661[129:66];
    assign _683 = PHASE_5 ? _682 : _681;
    assign _679 = _619[129:66];
    assign _678 = _605[129:66];
    assign q1_1 = PHASE_6 ? _679 : _678;
    assign _684 = _586 ? _683 : q1_1;
    assign address_26 = _663 ? _657 : _656;
    assign _669 = ~ _663;
    assign read_enable_20 = _102 & _669;
    assign address_27 = _663 ? _60 : _639;
    assign _665 = ~ _663;
    assign read_enable_21 = _102 & _665;
    assign _663 = ~ PHASE_5;
    assign write_enable_27 = _622 & _663;
    assign _667 = write_enable_27 | read_enable_21;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_12
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_667), .regcea(vdd), .wea(write_enable_27), .addra(address_27), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_20), .regceb(vdd), .web(write_enable_26), .addrb(address_26), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_674[131:131]), .sbiterrb(_674[130:130]), .doutb(_674[129:66]), .dbiterra(_674[65:65]), .sbiterra(_674[64:64]), .douta(_674[63:0]) );
    assign _675 = _674[63:0];
    assign _655 = _172[11:11];
    assign _654 = _172[10:10];
    assign _653 = _172[9:9];
    assign _652 = _172[8:8];
    assign _651 = _172[7:7];
    assign _650 = _172[6:6];
    assign _649 = _172[5:5];
    assign _648 = _172[4:4];
    assign _647 = _172[3:3];
    assign _646 = _172[2:2];
    assign _645 = _172[1:1];
    assign _644 = _172[0:0];
    assign _656 = { _644, _645, _646, _647, _648, _649, _650, _651, _652, _653, _654, _655 };
    assign address_28 = PHASE_5 ? _657 : _656;
    assign _641 = ~ PHASE_5;
    assign read_enable_22 = _102 & _641;
    assign data_25 = wr_d5;
    assign _638 = _137[11:11];
    assign _637 = _137[10:10];
    assign _636 = _137[9:9];
    assign _635 = _137[8:8];
    assign _634 = _137[7:7];
    assign _633 = _137[6:6];
    assign _632 = _137[5:5];
    assign _631 = _137[4:4];
    assign _630 = _137[3:3];
    assign _629 = _137[2:2];
    assign _628 = _137[1:1];
    assign _627 = _137[0:0];
    assign _639 = { _627, _628, _629, _630, _631, _632, _633, _634, _635, _636, _637, _638 };
    assign address_29 = PHASE_5 ? _60 : _639;
    assign _624 = ~ PHASE_5;
    assign read_enable_23 = _102 & _624;
    assign _622 = _62[5:5];
    assign write_enable_29 = _622 & PHASE_5;
    assign _626 = write_enable_29 | read_enable_23;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_13
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_626), .regcea(vdd), .wea(write_enable_29), .addra(address_29), .dina(data_25), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_22), .regceb(vdd), .web(write_enable_28), .addrb(address_28), .dinb(data_23), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_661[131:131]), .sbiterrb(_661[130:130]), .doutb(_661[129:66]), .dbiterra(_661[65:65]), .sbiterra(_661[64:64]), .douta(_661[63:0]) );
    assign _662 = _661[63:0];
    assign _583 = ~ PHASE_5;
    assign _19 = _583;
    always @(posedge _84) begin
        if (_82)
            PHASE_5 <= _581;
        else
            if (_72)
                PHASE_5 <= _19;
    end
    assign _676 = PHASE_5 ? _675 : _662;
    assign address_30 = _607 ? _199 : _172;
    assign _614 = ~ _607;
    assign read_enable_24 = _102 & _614;
    assign write_enable_30 = _598 & _607;
    assign _616 = write_enable_30 | read_enable_24;
    assign address_31 = _607 ? _164 : _137;
    assign _609 = ~ _607;
    assign read_enable_25 = _102 & _609;
    assign _607 = ~ PHASE_6;
    assign write_enable_31 = _591 & _607;
    assign _611 = write_enable_31 | read_enable_25;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_14
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_611), .regcea(vdd), .wea(write_enable_31), .addra(address_31), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_616), .regceb(vdd), .web(write_enable_30), .addrb(address_30), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_619[131:131]), .sbiterrb(_619[130:130]), .doutb(_619[129:66]), .dbiterra(_619[65:65]), .sbiterra(_619[64:64]), .douta(_619[63:0]) );
    assign _620 = _619[63:0];
    assign _687 = _686[127:64];
    assign data_27 = _687;
    assign address_32 = PHASE_6 ? _199 : _172;
    assign _600 = ~ PHASE_6;
    assign read_enable_26 = _102 & _600;
    assign _597 = ~ _130;
    assign _598 = _129 & _597;
    assign write_enable_32 = _598 & PHASE_6;
    assign _602 = write_enable_32 | read_enable_26;
    assign address_33 = PHASE_6 ? _164 : _137;
    assign _593 = ~ PHASE_6;
    assign read_enable_27 = _102 & _593;
    assign _590 = ~ _130;
    assign _591 = _129 & _590;
    assign write_enable_33 = _591 & PHASE_6;
    assign _595 = write_enable_33 | read_enable_27;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_15
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_595), .regcea(vdd), .wea(write_enable_33), .addra(address_33), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_602), .regceb(vdd), .web(write_enable_32), .addrb(address_32), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_605[131:131]), .sbiterrb(_605[130:130]), .doutb(_605[129:66]), .dbiterra(_605[65:65]), .sbiterra(_605[64:64]), .douta(_605[63:0]) );
    assign _606 = _605[63:0];
    assign _688 = ~ PHASE_6;
    assign _21 = _688;
    always @(posedge _84) begin
        if (_82)
            PHASE_6 <= _588;
        else
            if (_99)
                PHASE_6 <= _21;
    end
    assign q0_1 = PHASE_6 ? _620 : _606;
    always @(posedge _84) begin
        if (_82)
            _586 <= _585;
        else
            _586 <= _92;
    end
    assign _677 = _586 ? _676 : q0_1;
    dp_60
        dp_4
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_677), .d2(_684), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_686[191:128]), .q2(_686[127:64]), .q1(_686[63:0]) );
    assign _689 = _686[63:0];
    assign data_31 = _689;
    assign address_34 = PHASE_7 ? _164 : _68;
    assign _753 = ~ PHASE_7;
    assign _752 = _70[5:5];
    assign read_enable_28 = _752 & _753;
    always @(posedge _84) begin
        if (_82)
            _723 <= _722;
        else
            _723 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _726 <= _725;
        else
            _726 <= _723;
    end
    always @(posedge _84) begin
        if (_82)
            _729 <= _728;
        else
            _729 <= _726;
    end
    always @(posedge _84) begin
        if (_82)
            _732 <= _731;
        else
            _732 <= _729;
    end
    always @(posedge _84) begin
        if (_82)
            _735 <= _734;
        else
            _735 <= _732;
    end
    always @(posedge _84) begin
        if (_82)
            _738 <= _737;
        else
            _738 <= _735;
    end
    always @(posedge _84) begin
        if (_82)
            _741 <= _740;
        else
            _741 <= _738;
    end
    always @(posedge _84) begin
        if (_82)
            _744 <= _743;
        else
            _744 <= _741;
    end
    always @(posedge _84) begin
        if (_82)
            _747 <= _746;
        else
            _747 <= _744;
    end
    assign _748 = ~ _747;
    always @(posedge _84) begin
        if (_82)
            _696 <= _695;
        else
            _696 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _699 <= _698;
        else
            _699 <= _696;
    end
    always @(posedge _84) begin
        if (_82)
            _702 <= _701;
        else
            _702 <= _699;
    end
    always @(posedge _84) begin
        if (_82)
            _705 <= _704;
        else
            _705 <= _702;
    end
    always @(posedge _84) begin
        if (_82)
            _708 <= _707;
        else
            _708 <= _705;
    end
    always @(posedge _84) begin
        if (_82)
            _711 <= _710;
        else
            _711 <= _708;
    end
    always @(posedge _84) begin
        if (_82)
            _714 <= _713;
        else
            _714 <= _711;
    end
    always @(posedge _84) begin
        if (_82)
            _717 <= _716;
        else
            _717 <= _714;
    end
    always @(posedge _84) begin
        if (_82)
            _720 <= _719;
        else
            _720 <= _717;
    end
    assign _749 = _720 & _748;
    assign _750 = _129 & _749;
    assign write_enable_34 = _750 & PHASE_7;
    assign _755 = write_enable_34 | read_enable_28;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_16
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_755), .regcea(vdd), .wea(write_enable_34), .addra(address_34), .dina(data_31), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_25), .regceb(vdd), .web(write_enable_25), .addrb(address_25), .dinb(data_27), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_762[131:131]), .sbiterrb(_762[130:130]), .doutb(_762[129:66]), .dbiterra(_762[65:65]), .sbiterra(_762[64:64]), .douta(_762[63:0]) );
    assign _763 = _762[63:0];
    assign _693 = ~ PHASE_7;
    assign _23 = _693;
    always @(posedge _84) begin
        if (_82)
            PHASE_7 <= _691;
        else
            if (_72)
                PHASE_7 <= _23;
    end
    assign _775 = PHASE_7 ? _774 : _763;
    assign address_35 = _960 ? _199 : _955;
    assign write_enable_35 = _953 & _960;
    assign address_36 = _960 ? _164 : _68;
    assign _962 = ~ _960;
    assign read_enable_29 = _948 & _962;
    assign _960 = ~ PHASE_10;
    assign write_enable_36 = _946 & _960;
    assign _964 = write_enable_36 | read_enable_29;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_17
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_964), .regcea(vdd), .wea(write_enable_36), .addra(address_36), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_35), .regceb(vdd), .web(write_enable_35), .addrb(address_35), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_969[131:131]), .sbiterrb(_969[130:130]), .doutb(_969[129:66]), .dbiterra(_969[65:65]), .sbiterra(_969[64:64]), .douta(_969[63:0]) );
    assign _970 = _969[63:0];
    assign address_37 = PHASE_10 ? _199 : _955;
    assign _953 = _129 & _916;
    assign write_enable_37 = _953 & PHASE_10;
    assign _878 = _870[129:66];
    assign _877 = _857[129:66];
    assign _879 = PHASE_8 ? _878 : _877;
    assign _875 = _815[129:66];
    assign _874 = _801[129:66];
    assign q1_2 = PHASE_9 ? _875 : _874;
    assign _880 = _782 ? _879 : q1_2;
    assign address_38 = _859 ? _853 : _852;
    assign _865 = ~ _859;
    assign read_enable_30 = _102 & _865;
    assign address_39 = _859 ? _60 : _835;
    assign _861 = ~ _859;
    assign read_enable_31 = _102 & _861;
    assign _859 = ~ PHASE_8;
    assign write_enable_39 = _818 & _859;
    assign _863 = write_enable_39 | read_enable_31;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_18
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_863), .regcea(vdd), .wea(write_enable_39), .addra(address_39), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_30), .regceb(vdd), .web(write_enable_38), .addrb(address_38), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_870[131:131]), .sbiterrb(_870[130:130]), .doutb(_870[129:66]), .dbiterra(_870[65:65]), .sbiterra(_870[64:64]), .douta(_870[63:0]) );
    assign _871 = _870[63:0];
    assign _851 = _172[11:11];
    assign _850 = _172[10:10];
    assign _849 = _172[9:9];
    assign _848 = _172[8:8];
    assign _847 = _172[7:7];
    assign _846 = _172[6:6];
    assign _845 = _172[5:5];
    assign _844 = _172[4:4];
    assign _843 = _172[3:3];
    assign _842 = _172[2:2];
    assign _841 = _172[1:1];
    assign _840 = _172[0:0];
    assign _852 = { _840, _841, _842, _843, _844, _845, _846, _847, _848, _849, _850, _851 };
    assign address_40 = PHASE_8 ? _853 : _852;
    assign _837 = ~ PHASE_8;
    assign read_enable_32 = _102 & _837;
    assign data_37 = wr_d4;
    assign _834 = _137[11:11];
    assign _833 = _137[10:10];
    assign _832 = _137[9:9];
    assign _831 = _137[8:8];
    assign _830 = _137[7:7];
    assign _829 = _137[6:6];
    assign _828 = _137[5:5];
    assign _827 = _137[4:4];
    assign _826 = _137[3:3];
    assign _825 = _137[2:2];
    assign _824 = _137[1:1];
    assign _823 = _137[0:0];
    assign _835 = { _823, _824, _825, _826, _827, _828, _829, _830, _831, _832, _833, _834 };
    assign address_41 = PHASE_8 ? _60 : _835;
    assign _820 = ~ PHASE_8;
    assign read_enable_33 = _102 & _820;
    assign _818 = _62[4:4];
    assign write_enable_41 = _818 & PHASE_8;
    assign _822 = write_enable_41 | read_enable_33;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_19
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_822), .regcea(vdd), .wea(write_enable_41), .addra(address_41), .dina(data_37), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_32), .regceb(vdd), .web(write_enable_40), .addrb(address_40), .dinb(data_35), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_857[131:131]), .sbiterrb(_857[130:130]), .doutb(_857[129:66]), .dbiterra(_857[65:65]), .sbiterra(_857[64:64]), .douta(_857[63:0]) );
    assign _858 = _857[63:0];
    assign _779 = ~ PHASE_8;
    assign _27 = _779;
    always @(posedge _84) begin
        if (_82)
            PHASE_8 <= _777;
        else
            if (_72)
                PHASE_8 <= _27;
    end
    assign _872 = PHASE_8 ? _871 : _858;
    assign address_42 = _803 ? _199 : _172;
    assign _810 = ~ _803;
    assign read_enable_34 = _102 & _810;
    assign write_enable_42 = _794 & _803;
    assign _812 = write_enable_42 | read_enable_34;
    assign address_43 = _803 ? _164 : _137;
    assign _805 = ~ _803;
    assign read_enable_35 = _102 & _805;
    assign _803 = ~ PHASE_9;
    assign write_enable_43 = _787 & _803;
    assign _807 = write_enable_43 | read_enable_35;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_20
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_807), .regcea(vdd), .wea(write_enable_43), .addra(address_43), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_812), .regceb(vdd), .web(write_enable_42), .addrb(address_42), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_815[131:131]), .sbiterrb(_815[130:130]), .doutb(_815[129:66]), .dbiterra(_815[65:65]), .sbiterra(_815[64:64]), .douta(_815[63:0]) );
    assign _816 = _815[63:0];
    assign _883 = _882[127:64];
    assign data_39 = _883;
    assign address_44 = PHASE_9 ? _199 : _172;
    assign _796 = ~ PHASE_9;
    assign read_enable_36 = _102 & _796;
    assign _793 = ~ _130;
    assign _794 = _129 & _793;
    assign write_enable_44 = _794 & PHASE_9;
    assign _798 = write_enable_44 | read_enable_36;
    assign address_45 = PHASE_9 ? _164 : _137;
    assign _789 = ~ PHASE_9;
    assign read_enable_37 = _102 & _789;
    assign _786 = ~ _130;
    assign _787 = _129 & _786;
    assign write_enable_45 = _787 & PHASE_9;
    assign _791 = write_enable_45 | read_enable_37;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_21
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_791), .regcea(vdd), .wea(write_enable_45), .addra(address_45), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_798), .regceb(vdd), .web(write_enable_44), .addrb(address_44), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_801[131:131]), .sbiterrb(_801[130:130]), .doutb(_801[129:66]), .dbiterra(_801[65:65]), .sbiterra(_801[64:64]), .douta(_801[63:0]) );
    assign _802 = _801[63:0];
    assign _884 = ~ PHASE_9;
    assign _29 = _884;
    always @(posedge _84) begin
        if (_82)
            PHASE_9 <= _784;
        else
            if (_99)
                PHASE_9 <= _29;
    end
    assign q0_2 = PHASE_9 ? _816 : _802;
    always @(posedge _84) begin
        if (_82)
            _782 <= _781;
        else
            _782 <= _92;
    end
    assign _873 = _782 ? _872 : q0_2;
    dp_59
        dp_3
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_873), .d2(_880), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_882[191:128]), .q2(_882[127:64]), .q1(_882[63:0]) );
    assign _885 = _882[63:0];
    assign data_43 = _885;
    assign address_46 = PHASE_10 ? _164 : _68;
    assign _949 = ~ PHASE_10;
    assign _948 = _70[4:4];
    assign read_enable_38 = _948 & _949;
    always @(posedge _84) begin
        if (_82)
            _919 <= _918;
        else
            _919 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _922 <= _921;
        else
            _922 <= _919;
    end
    always @(posedge _84) begin
        if (_82)
            _925 <= _924;
        else
            _925 <= _922;
    end
    always @(posedge _84) begin
        if (_82)
            _928 <= _927;
        else
            _928 <= _925;
    end
    always @(posedge _84) begin
        if (_82)
            _931 <= _930;
        else
            _931 <= _928;
    end
    always @(posedge _84) begin
        if (_82)
            _934 <= _933;
        else
            _934 <= _931;
    end
    always @(posedge _84) begin
        if (_82)
            _937 <= _936;
        else
            _937 <= _934;
    end
    always @(posedge _84) begin
        if (_82)
            _940 <= _939;
        else
            _940 <= _937;
    end
    always @(posedge _84) begin
        if (_82)
            _943 <= _942;
        else
            _943 <= _940;
    end
    assign _944 = ~ _943;
    always @(posedge _84) begin
        if (_82)
            _892 <= _891;
        else
            _892 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _895 <= _894;
        else
            _895 <= _892;
    end
    always @(posedge _84) begin
        if (_82)
            _898 <= _897;
        else
            _898 <= _895;
    end
    always @(posedge _84) begin
        if (_82)
            _901 <= _900;
        else
            _901 <= _898;
    end
    always @(posedge _84) begin
        if (_82)
            _904 <= _903;
        else
            _904 <= _901;
    end
    always @(posedge _84) begin
        if (_82)
            _907 <= _906;
        else
            _907 <= _904;
    end
    always @(posedge _84) begin
        if (_82)
            _910 <= _909;
        else
            _910 <= _907;
    end
    always @(posedge _84) begin
        if (_82)
            _913 <= _912;
        else
            _913 <= _910;
    end
    always @(posedge _84) begin
        if (_82)
            _916 <= _915;
        else
            _916 <= _913;
    end
    assign _945 = _916 & _944;
    assign _946 = _129 & _945;
    assign write_enable_46 = _946 & PHASE_10;
    assign _951 = write_enable_46 | read_enable_38;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_22
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_951), .regcea(vdd), .wea(write_enable_46), .addra(address_46), .dina(data_43), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_37), .regceb(vdd), .web(write_enable_37), .addrb(address_37), .dinb(data_39), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_958[131:131]), .sbiterrb(_958[130:130]), .doutb(_958[129:66]), .dbiterra(_958[65:65]), .sbiterra(_958[64:64]), .douta(_958[63:0]) );
    assign _959 = _958[63:0];
    assign _889 = ~ PHASE_10;
    assign _31 = _889;
    always @(posedge _84) begin
        if (_82)
            PHASE_10 <= _887;
        else
            if (_72)
                PHASE_10 <= _31;
    end
    assign _971 = PHASE_10 ? _970 : _959;
    assign address_47 = _1156 ? _199 : _1151;
    assign write_enable_47 = _1149 & _1156;
    assign address_48 = _1156 ? _164 : _68;
    assign _1158 = ~ _1156;
    assign read_enable_39 = _1144 & _1158;
    assign _1156 = ~ PHASE_13;
    assign write_enable_48 = _1142 & _1156;
    assign _1160 = write_enable_48 | read_enable_39;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_23
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1160), .regcea(vdd), .wea(write_enable_48), .addra(address_48), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_47), .regceb(vdd), .web(write_enable_47), .addrb(address_47), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1165[131:131]), .sbiterrb(_1165[130:130]), .doutb(_1165[129:66]), .dbiterra(_1165[65:65]), .sbiterra(_1165[64:64]), .douta(_1165[63:0]) );
    assign _1166 = _1165[63:0];
    assign address_49 = PHASE_13 ? _199 : _1151;
    assign _1149 = _129 & _1112;
    assign write_enable_49 = _1149 & PHASE_13;
    assign _1074 = _1066[129:66];
    assign _1073 = _1053[129:66];
    assign _1075 = PHASE_11 ? _1074 : _1073;
    assign _1071 = _1011[129:66];
    assign _1070 = _997[129:66];
    assign q1_3 = PHASE_12 ? _1071 : _1070;
    assign _1076 = _978 ? _1075 : q1_3;
    assign address_50 = _1055 ? _1049 : _1048;
    assign _1061 = ~ _1055;
    assign read_enable_40 = _102 & _1061;
    assign address_51 = _1055 ? _60 : _1031;
    assign _1057 = ~ _1055;
    assign read_enable_41 = _102 & _1057;
    assign _1055 = ~ PHASE_11;
    assign write_enable_51 = _1014 & _1055;
    assign _1059 = write_enable_51 | read_enable_41;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_24
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1059), .regcea(vdd), .wea(write_enable_51), .addra(address_51), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_40), .regceb(vdd), .web(write_enable_50), .addrb(address_50), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1066[131:131]), .sbiterrb(_1066[130:130]), .doutb(_1066[129:66]), .dbiterra(_1066[65:65]), .sbiterra(_1066[64:64]), .douta(_1066[63:0]) );
    assign _1067 = _1066[63:0];
    assign _1047 = _172[11:11];
    assign _1046 = _172[10:10];
    assign _1045 = _172[9:9];
    assign _1044 = _172[8:8];
    assign _1043 = _172[7:7];
    assign _1042 = _172[6:6];
    assign _1041 = _172[5:5];
    assign _1040 = _172[4:4];
    assign _1039 = _172[3:3];
    assign _1038 = _172[2:2];
    assign _1037 = _172[1:1];
    assign _1036 = _172[0:0];
    assign _1048 = { _1036, _1037, _1038, _1039, _1040, _1041, _1042, _1043, _1044, _1045, _1046, _1047 };
    assign address_52 = PHASE_11 ? _1049 : _1048;
    assign _1033 = ~ PHASE_11;
    assign read_enable_42 = _102 & _1033;
    assign data_49 = wr_d3;
    assign _1030 = _137[11:11];
    assign _1029 = _137[10:10];
    assign _1028 = _137[9:9];
    assign _1027 = _137[8:8];
    assign _1026 = _137[7:7];
    assign _1025 = _137[6:6];
    assign _1024 = _137[5:5];
    assign _1023 = _137[4:4];
    assign _1022 = _137[3:3];
    assign _1021 = _137[2:2];
    assign _1020 = _137[1:1];
    assign _1019 = _137[0:0];
    assign _1031 = { _1019, _1020, _1021, _1022, _1023, _1024, _1025, _1026, _1027, _1028, _1029, _1030 };
    assign address_53 = PHASE_11 ? _60 : _1031;
    assign _1016 = ~ PHASE_11;
    assign read_enable_43 = _102 & _1016;
    assign _1014 = _62[3:3];
    assign write_enable_53 = _1014 & PHASE_11;
    assign _1018 = write_enable_53 | read_enable_43;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_25
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1018), .regcea(vdd), .wea(write_enable_53), .addra(address_53), .dina(data_49), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_42), .regceb(vdd), .web(write_enable_52), .addrb(address_52), .dinb(data_47), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1053[131:131]), .sbiterrb(_1053[130:130]), .doutb(_1053[129:66]), .dbiterra(_1053[65:65]), .sbiterra(_1053[64:64]), .douta(_1053[63:0]) );
    assign _1054 = _1053[63:0];
    assign _975 = ~ PHASE_11;
    assign _35 = _975;
    always @(posedge _84) begin
        if (_82)
            PHASE_11 <= _973;
        else
            if (_72)
                PHASE_11 <= _35;
    end
    assign _1068 = PHASE_11 ? _1067 : _1054;
    assign address_54 = _999 ? _199 : _172;
    assign _1006 = ~ _999;
    assign read_enable_44 = _102 & _1006;
    assign write_enable_54 = _990 & _999;
    assign _1008 = write_enable_54 | read_enable_44;
    assign address_55 = _999 ? _164 : _137;
    assign _1001 = ~ _999;
    assign read_enable_45 = _102 & _1001;
    assign _999 = ~ PHASE_12;
    assign write_enable_55 = _983 & _999;
    assign _1003 = write_enable_55 | read_enable_45;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_26
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1003), .regcea(vdd), .wea(write_enable_55), .addra(address_55), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1008), .regceb(vdd), .web(write_enable_54), .addrb(address_54), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1011[131:131]), .sbiterrb(_1011[130:130]), .doutb(_1011[129:66]), .dbiterra(_1011[65:65]), .sbiterra(_1011[64:64]), .douta(_1011[63:0]) );
    assign _1012 = _1011[63:0];
    assign _1079 = _1078[127:64];
    assign data_51 = _1079;
    assign address_56 = PHASE_12 ? _199 : _172;
    assign _992 = ~ PHASE_12;
    assign read_enable_46 = _102 & _992;
    assign _989 = ~ _130;
    assign _990 = _129 & _989;
    assign write_enable_56 = _990 & PHASE_12;
    assign _994 = write_enable_56 | read_enable_46;
    assign address_57 = PHASE_12 ? _164 : _137;
    assign _985 = ~ PHASE_12;
    assign read_enable_47 = _102 & _985;
    assign _982 = ~ _130;
    assign _983 = _129 & _982;
    assign write_enable_57 = _983 & PHASE_12;
    assign _987 = write_enable_57 | read_enable_47;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_27
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_987), .regcea(vdd), .wea(write_enable_57), .addra(address_57), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_994), .regceb(vdd), .web(write_enable_56), .addrb(address_56), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_997[131:131]), .sbiterrb(_997[130:130]), .doutb(_997[129:66]), .dbiterra(_997[65:65]), .sbiterra(_997[64:64]), .douta(_997[63:0]) );
    assign _998 = _997[63:0];
    assign _1080 = ~ PHASE_12;
    assign _37 = _1080;
    always @(posedge _84) begin
        if (_82)
            PHASE_12 <= _980;
        else
            if (_99)
                PHASE_12 <= _37;
    end
    assign q0_3 = PHASE_12 ? _1012 : _998;
    always @(posedge _84) begin
        if (_82)
            _978 <= _977;
        else
            _978 <= _92;
    end
    assign _1069 = _978 ? _1068 : q0_3;
    dp_58
        dp_2
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1069), .d2(_1076), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1078[191:128]), .q2(_1078[127:64]), .q1(_1078[63:0]) );
    assign _1081 = _1078[63:0];
    assign data_55 = _1081;
    assign address_58 = PHASE_13 ? _164 : _68;
    assign _1145 = ~ PHASE_13;
    assign _1144 = _70[3:3];
    assign read_enable_48 = _1144 & _1145;
    always @(posedge _84) begin
        if (_82)
            _1115 <= _1114;
        else
            _1115 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1118 <= _1117;
        else
            _1118 <= _1115;
    end
    always @(posedge _84) begin
        if (_82)
            _1121 <= _1120;
        else
            _1121 <= _1118;
    end
    always @(posedge _84) begin
        if (_82)
            _1124 <= _1123;
        else
            _1124 <= _1121;
    end
    always @(posedge _84) begin
        if (_82)
            _1127 <= _1126;
        else
            _1127 <= _1124;
    end
    always @(posedge _84) begin
        if (_82)
            _1130 <= _1129;
        else
            _1130 <= _1127;
    end
    always @(posedge _84) begin
        if (_82)
            _1133 <= _1132;
        else
            _1133 <= _1130;
    end
    always @(posedge _84) begin
        if (_82)
            _1136 <= _1135;
        else
            _1136 <= _1133;
    end
    always @(posedge _84) begin
        if (_82)
            _1139 <= _1138;
        else
            _1139 <= _1136;
    end
    assign _1140 = ~ _1139;
    always @(posedge _84) begin
        if (_82)
            _1088 <= _1087;
        else
            _1088 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1091 <= _1090;
        else
            _1091 <= _1088;
    end
    always @(posedge _84) begin
        if (_82)
            _1094 <= _1093;
        else
            _1094 <= _1091;
    end
    always @(posedge _84) begin
        if (_82)
            _1097 <= _1096;
        else
            _1097 <= _1094;
    end
    always @(posedge _84) begin
        if (_82)
            _1100 <= _1099;
        else
            _1100 <= _1097;
    end
    always @(posedge _84) begin
        if (_82)
            _1103 <= _1102;
        else
            _1103 <= _1100;
    end
    always @(posedge _84) begin
        if (_82)
            _1106 <= _1105;
        else
            _1106 <= _1103;
    end
    always @(posedge _84) begin
        if (_82)
            _1109 <= _1108;
        else
            _1109 <= _1106;
    end
    always @(posedge _84) begin
        if (_82)
            _1112 <= _1111;
        else
            _1112 <= _1109;
    end
    assign _1141 = _1112 & _1140;
    assign _1142 = _129 & _1141;
    assign write_enable_58 = _1142 & PHASE_13;
    assign _1147 = write_enable_58 | read_enable_48;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_28
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1147), .regcea(vdd), .wea(write_enable_58), .addra(address_58), .dina(data_55), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_49), .regceb(vdd), .web(write_enable_49), .addrb(address_49), .dinb(data_51), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1154[131:131]), .sbiterrb(_1154[130:130]), .doutb(_1154[129:66]), .dbiterra(_1154[65:65]), .sbiterra(_1154[64:64]), .douta(_1154[63:0]) );
    assign _1155 = _1154[63:0];
    assign _1085 = ~ PHASE_13;
    assign _39 = _1085;
    always @(posedge _84) begin
        if (_82)
            PHASE_13 <= _1083;
        else
            if (_72)
                PHASE_13 <= _39;
    end
    assign _1167 = PHASE_13 ? _1166 : _1155;
    assign address_59 = _1352 ? _199 : _1347;
    assign write_enable_59 = _1345 & _1352;
    assign address_60 = _1352 ? _164 : _68;
    assign _1354 = ~ _1352;
    assign read_enable_49 = _1340 & _1354;
    assign _1352 = ~ PHASE_16;
    assign write_enable_60 = _1338 & _1352;
    assign _1356 = write_enable_60 | read_enable_49;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_29
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1356), .regcea(vdd), .wea(write_enable_60), .addra(address_60), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_59), .regceb(vdd), .web(write_enable_59), .addrb(address_59), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1361[131:131]), .sbiterrb(_1361[130:130]), .doutb(_1361[129:66]), .dbiterra(_1361[65:65]), .sbiterra(_1361[64:64]), .douta(_1361[63:0]) );
    assign _1362 = _1361[63:0];
    assign address_61 = PHASE_16 ? _199 : _1347;
    assign _1345 = _129 & _1308;
    assign write_enable_61 = _1345 & PHASE_16;
    assign _1270 = _1262[129:66];
    assign _1269 = _1249[129:66];
    assign _1271 = PHASE_14 ? _1270 : _1269;
    assign _1267 = _1207[129:66];
    assign _1266 = _1193[129:66];
    assign q1_4 = PHASE_15 ? _1267 : _1266;
    assign _1272 = _1174 ? _1271 : q1_4;
    assign address_62 = _1251 ? _1245 : _1244;
    assign _1257 = ~ _1251;
    assign read_enable_50 = _102 & _1257;
    assign address_63 = _1251 ? _60 : _1227;
    assign _1253 = ~ _1251;
    assign read_enable_51 = _102 & _1253;
    assign _1251 = ~ PHASE_14;
    assign write_enable_63 = _1210 & _1251;
    assign _1255 = write_enable_63 | read_enable_51;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_30
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1255), .regcea(vdd), .wea(write_enable_63), .addra(address_63), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_50), .regceb(vdd), .web(write_enable_62), .addrb(address_62), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1262[131:131]), .sbiterrb(_1262[130:130]), .doutb(_1262[129:66]), .dbiterra(_1262[65:65]), .sbiterra(_1262[64:64]), .douta(_1262[63:0]) );
    assign _1263 = _1262[63:0];
    assign _1243 = _172[11:11];
    assign _1242 = _172[10:10];
    assign _1241 = _172[9:9];
    assign _1240 = _172[8:8];
    assign _1239 = _172[7:7];
    assign _1238 = _172[6:6];
    assign _1237 = _172[5:5];
    assign _1236 = _172[4:4];
    assign _1235 = _172[3:3];
    assign _1234 = _172[2:2];
    assign _1233 = _172[1:1];
    assign _1232 = _172[0:0];
    assign _1244 = { _1232, _1233, _1234, _1235, _1236, _1237, _1238, _1239, _1240, _1241, _1242, _1243 };
    assign address_64 = PHASE_14 ? _1245 : _1244;
    assign _1229 = ~ PHASE_14;
    assign read_enable_52 = _102 & _1229;
    assign data_61 = wr_d2;
    assign _1226 = _137[11:11];
    assign _1225 = _137[10:10];
    assign _1224 = _137[9:9];
    assign _1223 = _137[8:8];
    assign _1222 = _137[7:7];
    assign _1221 = _137[6:6];
    assign _1220 = _137[5:5];
    assign _1219 = _137[4:4];
    assign _1218 = _137[3:3];
    assign _1217 = _137[2:2];
    assign _1216 = _137[1:1];
    assign _1215 = _137[0:0];
    assign _1227 = { _1215, _1216, _1217, _1218, _1219, _1220, _1221, _1222, _1223, _1224, _1225, _1226 };
    assign address_65 = PHASE_14 ? _60 : _1227;
    assign _1212 = ~ PHASE_14;
    assign read_enable_53 = _102 & _1212;
    assign _1210 = _62[2:2];
    assign write_enable_65 = _1210 & PHASE_14;
    assign _1214 = write_enable_65 | read_enable_53;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_31
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1214), .regcea(vdd), .wea(write_enable_65), .addra(address_65), .dina(data_61), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_52), .regceb(vdd), .web(write_enable_64), .addrb(address_64), .dinb(data_59), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1249[131:131]), .sbiterrb(_1249[130:130]), .doutb(_1249[129:66]), .dbiterra(_1249[65:65]), .sbiterra(_1249[64:64]), .douta(_1249[63:0]) );
    assign _1250 = _1249[63:0];
    assign _1171 = ~ PHASE_14;
    assign _43 = _1171;
    always @(posedge _84) begin
        if (_82)
            PHASE_14 <= _1169;
        else
            if (_72)
                PHASE_14 <= _43;
    end
    assign _1264 = PHASE_14 ? _1263 : _1250;
    assign address_66 = _1195 ? _199 : _172;
    assign _1202 = ~ _1195;
    assign read_enable_54 = _102 & _1202;
    assign write_enable_66 = _1186 & _1195;
    assign _1204 = write_enable_66 | read_enable_54;
    assign address_67 = _1195 ? _164 : _137;
    assign _1197 = ~ _1195;
    assign read_enable_55 = _102 & _1197;
    assign _1195 = ~ PHASE_15;
    assign write_enable_67 = _1179 & _1195;
    assign _1199 = write_enable_67 | read_enable_55;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_32
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1199), .regcea(vdd), .wea(write_enable_67), .addra(address_67), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1204), .regceb(vdd), .web(write_enable_66), .addrb(address_66), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1207[131:131]), .sbiterrb(_1207[130:130]), .doutb(_1207[129:66]), .dbiterra(_1207[65:65]), .sbiterra(_1207[64:64]), .douta(_1207[63:0]) );
    assign _1208 = _1207[63:0];
    assign _1275 = _1274[127:64];
    assign data_63 = _1275;
    assign address_68 = PHASE_15 ? _199 : _172;
    assign _1188 = ~ PHASE_15;
    assign read_enable_56 = _102 & _1188;
    assign _1185 = ~ _130;
    assign _1186 = _129 & _1185;
    assign write_enable_68 = _1186 & PHASE_15;
    assign _1190 = write_enable_68 | read_enable_56;
    assign address_69 = PHASE_15 ? _164 : _137;
    assign _1181 = ~ PHASE_15;
    assign read_enable_57 = _102 & _1181;
    assign _1178 = ~ _130;
    assign _1179 = _129 & _1178;
    assign write_enable_69 = _1179 & PHASE_15;
    assign _1183 = write_enable_69 | read_enable_57;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_33
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1183), .regcea(vdd), .wea(write_enable_69), .addra(address_69), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1190), .regceb(vdd), .web(write_enable_68), .addrb(address_68), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1193[131:131]), .sbiterrb(_1193[130:130]), .doutb(_1193[129:66]), .dbiterra(_1193[65:65]), .sbiterra(_1193[64:64]), .douta(_1193[63:0]) );
    assign _1194 = _1193[63:0];
    assign _1276 = ~ PHASE_15;
    assign _45 = _1276;
    always @(posedge _84) begin
        if (_82)
            PHASE_15 <= _1176;
        else
            if (_99)
                PHASE_15 <= _45;
    end
    assign q0_4 = PHASE_15 ? _1208 : _1194;
    always @(posedge _84) begin
        if (_82)
            _1174 <= _1173;
        else
            _1174 <= _92;
    end
    assign _1265 = _1174 ? _1264 : q0_4;
    dp_57
        dp_1
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1265), .d2(_1272), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1274[191:128]), .q2(_1274[127:64]), .q1(_1274[63:0]) );
    assign _1277 = _1274[63:0];
    assign data_67 = _1277;
    assign address_70 = PHASE_16 ? _164 : _68;
    assign _1341 = ~ PHASE_16;
    assign _1340 = _70[2:2];
    assign read_enable_58 = _1340 & _1341;
    always @(posedge _84) begin
        if (_82)
            _1311 <= _1310;
        else
            _1311 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1314 <= _1313;
        else
            _1314 <= _1311;
    end
    always @(posedge _84) begin
        if (_82)
            _1317 <= _1316;
        else
            _1317 <= _1314;
    end
    always @(posedge _84) begin
        if (_82)
            _1320 <= _1319;
        else
            _1320 <= _1317;
    end
    always @(posedge _84) begin
        if (_82)
            _1323 <= _1322;
        else
            _1323 <= _1320;
    end
    always @(posedge _84) begin
        if (_82)
            _1326 <= _1325;
        else
            _1326 <= _1323;
    end
    always @(posedge _84) begin
        if (_82)
            _1329 <= _1328;
        else
            _1329 <= _1326;
    end
    always @(posedge _84) begin
        if (_82)
            _1332 <= _1331;
        else
            _1332 <= _1329;
    end
    always @(posedge _84) begin
        if (_82)
            _1335 <= _1334;
        else
            _1335 <= _1332;
    end
    assign _1336 = ~ _1335;
    always @(posedge _84) begin
        if (_82)
            _1284 <= _1283;
        else
            _1284 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1287 <= _1286;
        else
            _1287 <= _1284;
    end
    always @(posedge _84) begin
        if (_82)
            _1290 <= _1289;
        else
            _1290 <= _1287;
    end
    always @(posedge _84) begin
        if (_82)
            _1293 <= _1292;
        else
            _1293 <= _1290;
    end
    always @(posedge _84) begin
        if (_82)
            _1296 <= _1295;
        else
            _1296 <= _1293;
    end
    always @(posedge _84) begin
        if (_82)
            _1299 <= _1298;
        else
            _1299 <= _1296;
    end
    always @(posedge _84) begin
        if (_82)
            _1302 <= _1301;
        else
            _1302 <= _1299;
    end
    always @(posedge _84) begin
        if (_82)
            _1305 <= _1304;
        else
            _1305 <= _1302;
    end
    always @(posedge _84) begin
        if (_82)
            _1308 <= _1307;
        else
            _1308 <= _1305;
    end
    assign _1337 = _1308 & _1336;
    assign _1338 = _129 & _1337;
    assign write_enable_70 = _1338 & PHASE_16;
    assign _1343 = write_enable_70 | read_enable_58;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_34
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1343), .regcea(vdd), .wea(write_enable_70), .addra(address_70), .dina(data_67), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_61), .regceb(vdd), .web(write_enable_61), .addrb(address_61), .dinb(data_63), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1350[131:131]), .sbiterrb(_1350[130:130]), .doutb(_1350[129:66]), .dbiterra(_1350[65:65]), .sbiterra(_1350[64:64]), .douta(_1350[63:0]) );
    assign _1351 = _1350[63:0];
    assign _1281 = ~ PHASE_16;
    assign _47 = _1281;
    always @(posedge _84) begin
        if (_82)
            PHASE_16 <= _1279;
        else
            if (_72)
                PHASE_16 <= _47;
    end
    assign _1363 = PHASE_16 ? _1362 : _1351;
    assign address_71 = _1548 ? _199 : _1543;
    assign write_enable_71 = _1541 & _1548;
    assign address_72 = _1548 ? _164 : _68;
    assign _1550 = ~ _1548;
    assign read_enable_59 = _1536 & _1550;
    assign _1548 = ~ PHASE_19;
    assign write_enable_72 = _1534 & _1548;
    assign _1552 = write_enable_72 | read_enable_59;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_35
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1552), .regcea(vdd), .wea(write_enable_72), .addra(address_72), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_71), .regceb(vdd), .web(write_enable_71), .addrb(address_71), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1557[131:131]), .sbiterrb(_1557[130:130]), .doutb(_1557[129:66]), .dbiterra(_1557[65:65]), .sbiterra(_1557[64:64]), .douta(_1557[63:0]) );
    assign _1558 = _1557[63:0];
    assign address_73 = PHASE_19 ? _199 : _1543;
    assign _1541 = _129 & _1504;
    assign write_enable_73 = _1541 & PHASE_19;
    assign _1466 = _1458[129:66];
    assign _1465 = _1445[129:66];
    assign _1467 = PHASE_17 ? _1466 : _1465;
    assign _1463 = _1403[129:66];
    assign _1462 = _1389[129:66];
    assign q1_5 = PHASE_18 ? _1463 : _1462;
    assign _1468 = _1370 ? _1467 : q1_5;
    assign address_74 = _1447 ? _1441 : _1440;
    assign _1453 = ~ _1447;
    assign read_enable_60 = _102 & _1453;
    assign address_75 = _1447 ? _60 : _1423;
    assign _1449 = ~ _1447;
    assign read_enable_61 = _102 & _1449;
    assign _1447 = ~ PHASE_17;
    assign write_enable_75 = _1406 & _1447;
    assign _1451 = write_enable_75 | read_enable_61;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_36
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1451), .regcea(vdd), .wea(write_enable_75), .addra(address_75), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_60), .regceb(vdd), .web(write_enable_74), .addrb(address_74), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1458[131:131]), .sbiterrb(_1458[130:130]), .doutb(_1458[129:66]), .dbiterra(_1458[65:65]), .sbiterra(_1458[64:64]), .douta(_1458[63:0]) );
    assign _1459 = _1458[63:0];
    assign _1439 = _172[11:11];
    assign _1438 = _172[10:10];
    assign _1437 = _172[9:9];
    assign _1436 = _172[8:8];
    assign _1435 = _172[7:7];
    assign _1434 = _172[6:6];
    assign _1433 = _172[5:5];
    assign _1432 = _172[4:4];
    assign _1431 = _172[3:3];
    assign _1430 = _172[2:2];
    assign _1429 = _172[1:1];
    assign _1428 = _172[0:0];
    assign _1440 = { _1428, _1429, _1430, _1431, _1432, _1433, _1434, _1435, _1436, _1437, _1438, _1439 };
    assign address_76 = PHASE_17 ? _1441 : _1440;
    assign _1425 = ~ PHASE_17;
    assign read_enable_62 = _102 & _1425;
    assign data_73 = wr_d1;
    assign _1422 = _137[11:11];
    assign _1421 = _137[10:10];
    assign _1420 = _137[9:9];
    assign _1419 = _137[8:8];
    assign _1418 = _137[7:7];
    assign _1417 = _137[6:6];
    assign _1416 = _137[5:5];
    assign _1415 = _137[4:4];
    assign _1414 = _137[3:3];
    assign _1413 = _137[2:2];
    assign _1412 = _137[1:1];
    assign _1411 = _137[0:0];
    assign _1423 = { _1411, _1412, _1413, _1414, _1415, _1416, _1417, _1418, _1419, _1420, _1421, _1422 };
    assign address_77 = PHASE_17 ? _60 : _1423;
    assign _1408 = ~ PHASE_17;
    assign read_enable_63 = _102 & _1408;
    assign _1406 = _62[1:1];
    assign write_enable_77 = _1406 & PHASE_17;
    assign _1410 = write_enable_77 | read_enable_63;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_37
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1410), .regcea(vdd), .wea(write_enable_77), .addra(address_77), .dina(data_73), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_62), .regceb(vdd), .web(write_enable_76), .addrb(address_76), .dinb(data_71), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1445[131:131]), .sbiterrb(_1445[130:130]), .doutb(_1445[129:66]), .dbiterra(_1445[65:65]), .sbiterra(_1445[64:64]), .douta(_1445[63:0]) );
    assign _1446 = _1445[63:0];
    assign _1367 = ~ PHASE_17;
    assign _51 = _1367;
    always @(posedge _84) begin
        if (_82)
            PHASE_17 <= _1365;
        else
            if (_72)
                PHASE_17 <= _51;
    end
    assign _1460 = PHASE_17 ? _1459 : _1446;
    assign address_78 = _1391 ? _199 : _172;
    assign _1398 = ~ _1391;
    assign read_enable_64 = _102 & _1398;
    assign write_enable_78 = _1382 & _1391;
    assign _1400 = write_enable_78 | read_enable_64;
    assign address_79 = _1391 ? _164 : _137;
    assign _1393 = ~ _1391;
    assign read_enable_65 = _102 & _1393;
    assign _1391 = ~ PHASE_18;
    assign write_enable_79 = _1375 & _1391;
    assign _1395 = write_enable_79 | read_enable_65;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_38
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1395), .regcea(vdd), .wea(write_enable_79), .addra(address_79), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1400), .regceb(vdd), .web(write_enable_78), .addrb(address_78), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1403[131:131]), .sbiterrb(_1403[130:130]), .doutb(_1403[129:66]), .dbiterra(_1403[65:65]), .sbiterra(_1403[64:64]), .douta(_1403[63:0]) );
    assign _1404 = _1403[63:0];
    assign _1471 = _1470[127:64];
    assign data_75 = _1471;
    assign address_80 = PHASE_18 ? _199 : _172;
    assign _1384 = ~ PHASE_18;
    assign read_enable_66 = _102 & _1384;
    assign _1381 = ~ _130;
    assign _1382 = _129 & _1381;
    assign write_enable_80 = _1382 & PHASE_18;
    assign _1386 = write_enable_80 | read_enable_66;
    assign address_81 = PHASE_18 ? _164 : _137;
    assign _1377 = ~ PHASE_18;
    assign read_enable_67 = _102 & _1377;
    assign _1374 = ~ _130;
    assign _1375 = _129 & _1374;
    assign write_enable_81 = _1375 & PHASE_18;
    assign _1379 = write_enable_81 | read_enable_67;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_39
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1379), .regcea(vdd), .wea(write_enable_81), .addra(address_81), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1386), .regceb(vdd), .web(write_enable_80), .addrb(address_80), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1389[131:131]), .sbiterrb(_1389[130:130]), .doutb(_1389[129:66]), .dbiterra(_1389[65:65]), .sbiterra(_1389[64:64]), .douta(_1389[63:0]) );
    assign _1390 = _1389[63:0];
    assign _1472 = ~ PHASE_18;
    assign _53 = _1472;
    always @(posedge _84) begin
        if (_82)
            PHASE_18 <= _1372;
        else
            if (_99)
                PHASE_18 <= _53;
    end
    assign q0_5 = PHASE_18 ? _1404 : _1390;
    always @(posedge _84) begin
        if (_82)
            _1370 <= _1369;
        else
            _1370 <= _92;
    end
    assign _1461 = _1370 ? _1460 : q0_5;
    dp_56
        dp_0
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1461), .d2(_1468), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1470[191:128]), .q2(_1470[127:64]), .q1(_1470[63:0]) );
    assign _1473 = _1470[63:0];
    assign data_79 = _1473;
    assign address_82 = PHASE_19 ? _164 : _68;
    assign _1537 = ~ PHASE_19;
    assign _1536 = _70[1:1];
    assign read_enable_68 = _1536 & _1537;
    always @(posedge _84) begin
        if (_82)
            _1507 <= _1506;
        else
            _1507 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1510 <= _1509;
        else
            _1510 <= _1507;
    end
    always @(posedge _84) begin
        if (_82)
            _1513 <= _1512;
        else
            _1513 <= _1510;
    end
    always @(posedge _84) begin
        if (_82)
            _1516 <= _1515;
        else
            _1516 <= _1513;
    end
    always @(posedge _84) begin
        if (_82)
            _1519 <= _1518;
        else
            _1519 <= _1516;
    end
    always @(posedge _84) begin
        if (_82)
            _1522 <= _1521;
        else
            _1522 <= _1519;
    end
    always @(posedge _84) begin
        if (_82)
            _1525 <= _1524;
        else
            _1525 <= _1522;
    end
    always @(posedge _84) begin
        if (_82)
            _1528 <= _1527;
        else
            _1528 <= _1525;
    end
    always @(posedge _84) begin
        if (_82)
            _1531 <= _1530;
        else
            _1531 <= _1528;
    end
    assign _1532 = ~ _1531;
    always @(posedge _84) begin
        if (_82)
            _1480 <= _1479;
        else
            _1480 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1483 <= _1482;
        else
            _1483 <= _1480;
    end
    always @(posedge _84) begin
        if (_82)
            _1486 <= _1485;
        else
            _1486 <= _1483;
    end
    always @(posedge _84) begin
        if (_82)
            _1489 <= _1488;
        else
            _1489 <= _1486;
    end
    always @(posedge _84) begin
        if (_82)
            _1492 <= _1491;
        else
            _1492 <= _1489;
    end
    always @(posedge _84) begin
        if (_82)
            _1495 <= _1494;
        else
            _1495 <= _1492;
    end
    always @(posedge _84) begin
        if (_82)
            _1498 <= _1497;
        else
            _1498 <= _1495;
    end
    always @(posedge _84) begin
        if (_82)
            _1501 <= _1500;
        else
            _1501 <= _1498;
    end
    always @(posedge _84) begin
        if (_82)
            _1504 <= _1503;
        else
            _1504 <= _1501;
    end
    assign _1533 = _1504 & _1532;
    assign _1534 = _129 & _1533;
    assign write_enable_82 = _1534 & PHASE_19;
    assign _1539 = write_enable_82 | read_enable_68;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_40
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1539), .regcea(vdd), .wea(write_enable_82), .addra(address_82), .dina(data_79), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_73), .regceb(vdd), .web(write_enable_73), .addrb(address_73), .dinb(data_75), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1546[131:131]), .sbiterrb(_1546[130:130]), .doutb(_1546[129:66]), .dbiterra(_1546[65:65]), .sbiterra(_1546[64:64]), .douta(_1546[63:0]) );
    assign _1547 = _1546[63:0];
    assign _1477 = ~ PHASE_19;
    assign _55 = _1477;
    always @(posedge _84) begin
        if (_82)
            PHASE_19 <= _1475;
        else
            if (_72)
                PHASE_19 <= _55;
    end
    assign _1559 = PHASE_19 ? _1558 : _1547;
    assign address_83 = _1744 ? _199 : _1739;
    assign write_enable_83 = _1737 & _1744;
    assign address_84 = _1744 ? _164 : _68;
    assign _1746 = ~ _1744;
    assign read_enable_69 = _1732 & _1746;
    assign _1744 = ~ PHASE_22;
    assign write_enable_84 = _1730 & _1744;
    assign _1748 = write_enable_84 | read_enable_69;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_41
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1748), .regcea(vdd), .wea(write_enable_84), .addra(address_84), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_83), .regceb(vdd), .web(write_enable_83), .addrb(address_83), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1753[131:131]), .sbiterrb(_1753[130:130]), .doutb(_1753[129:66]), .dbiterra(_1753[65:65]), .sbiterra(_1753[64:64]), .douta(_1753[63:0]) );
    assign _1754 = _1753[63:0];
    assign address_85 = PHASE_22 ? _199 : _1739;
    assign _1737 = _129 & _1700;
    assign write_enable_85 = _1737 & PHASE_22;
    assign _292 = _91[521:518];
    assign _291 = _91[517:517];
    assign _289 = _91[513:513];
    assign _288 = _91[512:449];
    assign _287 = _91[448:385];
    assign _286 = _91[384:321];
    assign _285 = _91[320:257];
    assign _284 = _91[256:193];
    assign _283 = _91[192:129];
    assign _282 = _91[128:65];
    assign _1662 = _1654[129:66];
    assign _1661 = _1641[129:66];
    assign _1663 = PHASE_20 ? _1662 : _1661;
    assign _1659 = _1599[129:66];
    assign _1658 = _1585[129:66];
    assign q1_6 = PHASE_21 ? _1659 : _1658;
    assign _1664 = _1566 ? _1663 : q1_6;
    assign address_86 = _1643 ? _1637 : _1636;
    assign _1649 = ~ _1643;
    assign read_enable_70 = _102 & _1649;
    assign address_87 = _1643 ? _60 : _1619;
    assign _1645 = ~ _1643;
    assign read_enable_71 = _102 & _1645;
    assign _1643 = ~ PHASE_20;
    assign write_enable_87 = _1602 & _1643;
    assign _1647 = write_enable_87 | read_enable_71;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_42
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1647), .regcea(vdd), .wea(write_enable_87), .addra(address_87), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_70), .regceb(vdd), .web(write_enable_86), .addrb(address_86), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1654[131:131]), .sbiterrb(_1654[130:130]), .doutb(_1654[129:66]), .dbiterra(_1654[65:65]), .sbiterra(_1654[64:64]), .douta(_1654[63:0]) );
    assign _1655 = _1654[63:0];
    assign _1635 = _172[11:11];
    assign _1634 = _172[10:10];
    assign _1633 = _172[9:9];
    assign _1632 = _172[8:8];
    assign _1631 = _172[7:7];
    assign _1630 = _172[6:6];
    assign _1629 = _172[5:5];
    assign _1628 = _172[4:4];
    assign _1627 = _172[3:3];
    assign _1626 = _172[2:2];
    assign _1625 = _172[1:1];
    assign _1624 = _172[0:0];
    assign _1636 = { _1624, _1625, _1626, _1627, _1628, _1629, _1630, _1631, _1632, _1633, _1634, _1635 };
    assign address_88 = PHASE_20 ? _1637 : _1636;
    assign _1621 = ~ PHASE_20;
    assign read_enable_72 = _102 & _1621;
    assign data_85 = wr_d0;
    assign _60 = wr_addr;
    assign _1618 = _137[11:11];
    assign _1617 = _137[10:10];
    assign _1616 = _137[9:9];
    assign _1615 = _137[8:8];
    assign _1614 = _137[7:7];
    assign _1613 = _137[6:6];
    assign _1612 = _137[5:5];
    assign _1611 = _137[4:4];
    assign _1610 = _137[3:3];
    assign _1609 = _137[2:2];
    assign _1608 = _137[1:1];
    assign _1607 = _137[0:0];
    assign _1619 = { _1607, _1608, _1609, _1610, _1611, _1612, _1613, _1614, _1615, _1616, _1617, _1618 };
    assign address_89 = PHASE_20 ? _60 : _1619;
    assign _1604 = ~ PHASE_20;
    assign read_enable_73 = _102 & _1604;
    assign _62 = wr_en;
    assign _1602 = _62[0:0];
    assign write_enable_89 = _1602 & PHASE_20;
    assign _1606 = write_enable_89 | read_enable_73;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_43
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1606), .regcea(vdd), .wea(write_enable_89), .addra(address_89), .dina(data_85), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(read_enable_72), .regceb(vdd), .web(write_enable_88), .addrb(address_88), .dinb(data_83), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1641[131:131]), .sbiterrb(_1641[130:130]), .doutb(_1641[129:66]), .dbiterra(_1641[65:65]), .sbiterra(_1641[64:64]), .douta(_1641[63:0]) );
    assign _1642 = _1641[63:0];
    assign _1563 = ~ PHASE_20;
    assign _63 = _1563;
    always @(posedge _84) begin
        if (_82)
            PHASE_20 <= _1561;
        else
            if (_72)
                PHASE_20 <= _63;
    end
    assign _1656 = PHASE_20 ? _1655 : _1642;
    assign address_90 = _1587 ? _199 : _172;
    assign _1594 = ~ _1587;
    assign read_enable_74 = _102 & _1594;
    assign write_enable_90 = _1578 & _1587;
    assign _1596 = write_enable_90 | read_enable_74;
    assign address_91 = _1587 ? _164 : _137;
    assign _1589 = ~ _1587;
    assign read_enable_75 = _102 & _1589;
    assign _1587 = ~ PHASE_21;
    assign write_enable_91 = _1571 & _1587;
    assign _1591 = write_enable_91 | read_enable_75;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_44
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1591), .regcea(vdd), .wea(write_enable_91), .addra(address_91), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1596), .regceb(vdd), .web(write_enable_90), .addrb(address_90), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1599[131:131]), .sbiterrb(_1599[130:130]), .doutb(_1599[129:66]), .dbiterra(_1599[65:65]), .sbiterra(_1599[64:64]), .douta(_1599[63:0]) );
    assign _1600 = _1599[63:0];
    assign _1667 = _1666[127:64];
    assign data_87 = _1667;
    always @(posedge _84) begin
        if (_82)
            _175 <= _174;
        else
            _175 <= _172;
    end
    always @(posedge _84) begin
        if (_82)
            _178 <= _177;
        else
            _178 <= _175;
    end
    always @(posedge _84) begin
        if (_82)
            _181 <= _180;
        else
            _181 <= _178;
    end
    always @(posedge _84) begin
        if (_82)
            _184 <= _183;
        else
            _184 <= _181;
    end
    always @(posedge _84) begin
        if (_82)
            _187 <= _186;
        else
            _187 <= _184;
    end
    always @(posedge _84) begin
        if (_82)
            _190 <= _189;
        else
            _190 <= _187;
    end
    always @(posedge _84) begin
        if (_82)
            _193 <= _192;
        else
            _193 <= _190;
    end
    always @(posedge _84) begin
        if (_82)
            _196 <= _195;
        else
            _196 <= _193;
    end
    always @(posedge _84) begin
        if (_82)
            _199 <= _198;
        else
            _199 <= _196;
    end
    assign _172 = _91[64:53];
    assign address_92 = PHASE_21 ? _199 : _172;
    assign _1580 = ~ PHASE_21;
    assign read_enable_76 = _102 & _1580;
    assign _1577 = ~ _130;
    assign _1578 = _129 & _1577;
    assign write_enable_92 = _1578 & PHASE_21;
    assign _1582 = write_enable_92 | read_enable_76;
    assign address_93 = PHASE_21 ? _164 : _137;
    assign _1573 = ~ PHASE_21;
    assign read_enable_77 = _102 & _1573;
    assign _1570 = ~ _130;
    assign _1571 = _129 & _1570;
    assign write_enable_93 = _1571 & PHASE_21;
    assign _1575 = write_enable_93 | read_enable_77;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_45
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1575), .regcea(vdd), .wea(write_enable_93), .addra(address_93), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(_1582), .regceb(vdd), .web(write_enable_92), .addrb(address_92), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1585[131:131]), .sbiterrb(_1585[130:130]), .doutb(_1585[129:66]), .dbiterra(_1585[65:65]), .sbiterra(_1585[64:64]), .douta(_1585[63:0]) );
    assign _1586 = _1585[63:0];
    assign _99 = _91[523:523];
    assign _1668 = ~ PHASE_21;
    assign _65 = _1668;
    always @(posedge _84) begin
        if (_82)
            PHASE_21 <= _1568;
        else
            if (_99)
                PHASE_21 <= _65;
    end
    assign q0_6 = PHASE_21 ? _1600 : _1586;
    assign _92 = _91[514:514];
    always @(posedge _84) begin
        if (_82)
            _1566 <= _1565;
        else
            _1566 <= _92;
    end
    assign _1657 = _1566 ? _1656 : q0_6;
    dp_55
        dp
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .d1(_1657), .d2(_1664), .omegas0(_282), .omegas1(_283), .omegas2(_284), .omegas3(_285), .omegas4(_286), .omegas5(_287), .omegas6(_288), .start_twiddles(_289), .twiddle_stage(_290), .valid(_291), .index(_292), .twiddle_update_q(_1666[191:128]), .q2(_1666[127:64]), .q1(_1666[63:0]) );
    assign _1669 = _1666[63:0];
    assign data_91 = _1669;
    assign _137 = _91[52:41];
    always @(posedge _84) begin
        if (_82)
            _140 <= _139;
        else
            _140 <= _137;
    end
    always @(posedge _84) begin
        if (_82)
            _143 <= _142;
        else
            _143 <= _140;
    end
    always @(posedge _84) begin
        if (_82)
            _146 <= _145;
        else
            _146 <= _143;
    end
    always @(posedge _84) begin
        if (_82)
            _149 <= _148;
        else
            _149 <= _146;
    end
    always @(posedge _84) begin
        if (_82)
            _152 <= _151;
        else
            _152 <= _149;
    end
    always @(posedge _84) begin
        if (_82)
            _155 <= _154;
        else
            _155 <= _152;
    end
    always @(posedge _84) begin
        if (_82)
            _158 <= _157;
        else
            _158 <= _155;
    end
    always @(posedge _84) begin
        if (_82)
            _161 <= _160;
        else
            _161 <= _158;
    end
    always @(posedge _84) begin
        if (_82)
            _164 <= _163;
        else
            _164 <= _161;
    end
    assign _68 = rd_addr;
    assign address_94 = PHASE_22 ? _164 : _68;
    assign _1733 = ~ PHASE_22;
    assign _70 = rd_en;
    assign _1732 = _70[0:0];
    assign read_enable_78 = _1732 & _1733;
    assign _290 = _91[516:516];
    always @(posedge _84) begin
        if (_82)
            _1703 <= _1702;
        else
            _1703 <= _290;
    end
    always @(posedge _84) begin
        if (_82)
            _1706 <= _1705;
        else
            _1706 <= _1703;
    end
    always @(posedge _84) begin
        if (_82)
            _1709 <= _1708;
        else
            _1709 <= _1706;
    end
    always @(posedge _84) begin
        if (_82)
            _1712 <= _1711;
        else
            _1712 <= _1709;
    end
    always @(posedge _84) begin
        if (_82)
            _1715 <= _1714;
        else
            _1715 <= _1712;
    end
    always @(posedge _84) begin
        if (_82)
            _1718 <= _1717;
        else
            _1718 <= _1715;
    end
    always @(posedge _84) begin
        if (_82)
            _1721 <= _1720;
        else
            _1721 <= _1718;
    end
    always @(posedge _84) begin
        if (_82)
            _1724 <= _1723;
        else
            _1724 <= _1721;
    end
    always @(posedge _84) begin
        if (_82)
            _1727 <= _1726;
        else
            _1727 <= _1724;
    end
    assign _1728 = ~ _1727;
    assign _130 = _91[515:515];
    always @(posedge _84) begin
        if (_82)
            _1676 <= _1675;
        else
            _1676 <= _130;
    end
    always @(posedge _84) begin
        if (_82)
            _1679 <= _1678;
        else
            _1679 <= _1676;
    end
    always @(posedge _84) begin
        if (_82)
            _1682 <= _1681;
        else
            _1682 <= _1679;
    end
    always @(posedge _84) begin
        if (_82)
            _1685 <= _1684;
        else
            _1685 <= _1682;
    end
    always @(posedge _84) begin
        if (_82)
            _1688 <= _1687;
        else
            _1688 <= _1685;
    end
    always @(posedge _84) begin
        if (_82)
            _1691 <= _1690;
        else
            _1691 <= _1688;
    end
    always @(posedge _84) begin
        if (_82)
            _1694 <= _1693;
        else
            _1694 <= _1691;
    end
    always @(posedge _84) begin
        if (_82)
            _1697 <= _1696;
        else
            _1697 <= _1694;
    end
    always @(posedge _84) begin
        if (_82)
            _1700 <= _1699;
        else
            _1700 <= _1697;
    end
    assign _1729 = _1700 & _1728;
    assign _102 = _91[522:522];
    always @(posedge _84) begin
        if (_82)
            _105 <= _104;
        else
            _105 <= _102;
    end
    always @(posedge _84) begin
        if (_82)
            _108 <= _107;
        else
            _108 <= _105;
    end
    always @(posedge _84) begin
        if (_82)
            _111 <= _110;
        else
            _111 <= _108;
    end
    always @(posedge _84) begin
        if (_82)
            _114 <= _113;
        else
            _114 <= _111;
    end
    always @(posedge _84) begin
        if (_82)
            _117 <= _116;
        else
            _117 <= _114;
    end
    always @(posedge _84) begin
        if (_82)
            _120 <= _119;
        else
            _120 <= _117;
    end
    always @(posedge _84) begin
        if (_82)
            _123 <= _122;
        else
            _123 <= _120;
    end
    always @(posedge _84) begin
        if (_82)
            _126 <= _125;
        else
            _126 <= _123;
    end
    always @(posedge _84) begin
        if (_82)
            _129 <= _128;
        else
            _129 <= _126;
    end
    assign _1730 = _129 & _1729;
    assign write_enable_94 = _1730 & PHASE_22;
    assign _1735 = write_enable_94 | read_enable_78;
    xpm_memory_tdpram
        #( .MEMORY_SIZE(262144), .MEMORY_PRIMITIVE("ultra"), .CLOCKING_MODE("common_clock"), .ECC_MODE("no_ecc"), .MEMORY_INIT_FILE("none"), .MEMORY_INIT_PARAM(""), .USE_MEM_INIT(0), .WAKEUP_TIME("disable_sleep"), .AUTO_SLEEP_TIME(0), .MESSAGE_CONTROL(0), .USE_EMBEDDED_CONSTRAINT(0), .MEMORY_OPTIMIZATION("true"), .CASCADE_HEIGHT(0), .SIM_ASSERT_CHK(0), .WRITE_DATA_WIDTH_A(64), .READ_DATA_WIDTH_A(64), .BYTE_WRITE_WIDTH_A(64), .ADDR_WIDTH_A(12), .READ_RESET_VALUE_A("0"), .READ_LATENCY_A(1), .WRITE_MODE_A("no_change"), .RST_MODE_A("SYNC"), .WRITE_DATA_WIDTH_B(64), .READ_DATA_WIDTH_B(64), .BYTE_WRITE_WIDTH_B(64), .ADDR_WIDTH_B(12), .READ_RESET_VALUE_B("0"), .READ_LATENCY_B(1), .WRITE_MODE_B("no_change"), .RST_MODE_B("SYNC") )
        the_xpm_memory_tdpram_46
        ( .sleep(gnd), .clka(_84), .rsta(gnd), .ena(_1735), .regcea(vdd), .wea(write_enable_94), .addra(address_94), .dina(data_91), .injectsbiterra(gnd), .injectdbiterra(gnd), .clkb(_84), .rstb(gnd), .enb(write_enable_85), .regceb(vdd), .web(write_enable_85), .addrb(address_85), .dinb(data_87), .injectsbiterrb(gnd), .injectdbiterrb(gnd), .dbiterrb(_1742[131:131]), .sbiterrb(_1742[130:130]), .doutb(_1742[129:66]), .dbiterra(_1742[65:65]), .sbiterra(_1742[64:64]), .douta(_1742[63:0]) );
    assign _1743 = _1742[63:0];
    assign _72 = flip;
    assign _1673 = ~ PHASE_22;
    assign _73 = _1673;
    always @(posedge _84) begin
        if (_82)
            PHASE_22 <= _1671;
        else
            if (_72)
                PHASE_22 <= _73;
    end
    assign _1755 = PHASE_22 ? _1754 : _1743;
    assign _76 = first_4step_pass;
    assign _78 = first_iter;
    assign _80 = start;
    assign _82 = clear;
    assign _84 = clock;
    ctrl
        ctrl
        ( .clock(_84), .clear(_82), .start(_80), .first_iter(_78), .first_4step_pass(_76), .flip(_91[523:523]), .read_write_enable(_91[522:522]), .index(_91[521:518]), .valid(_91[517:517]), .twiddle_stage(_91[516:516]), .last_stage(_91[515:515]), .first_stage(_91[514:514]), .start_twiddles(_91[513:513]), .omegas6(_91[512:449]), .omegas5(_91[448:385]), .omegas4(_91[384:321]), .omegas3(_91[320:257]), .omegas2(_91[256:193]), .omegas1(_91[192:129]), .omegas0(_91[128:65]), .addr2(_91[64:53]), .addr1(_91[52:41]), .m(_91[40:29]), .k(_91[28:17]), .j(_91[16:5]), .i(_91[4:1]), .done_(_91[0:0]) );
    assign _1756 = _91[0:0];

    /* aliases */
    assign data_0 = data;
    assign data_2 = data_1;
    assign data_4 = data_3;
    assign data_5 = data_3;
    assign data_6 = data_3;
    assign data_8 = data_7;
    assign data_9 = data_7;
    assign data_10 = data_7;
    assign data_12 = data_11;
    assign data_14 = data_13;
    assign data_16 = data_15;
    assign data_17 = data_15;
    assign data_18 = data_15;
    assign data_20 = data_19;
    assign data_21 = data_19;
    assign data_22 = data_19;
    assign data_24 = data_23;
    assign data_26 = data_25;
    assign data_28 = data_27;
    assign data_29 = data_27;
    assign data_30 = data_27;
    assign data_32 = data_31;
    assign data_33 = data_31;
    assign data_34 = data_31;
    assign data_36 = data_35;
    assign data_38 = data_37;
    assign data_40 = data_39;
    assign data_41 = data_39;
    assign data_42 = data_39;
    assign data_44 = data_43;
    assign data_45 = data_43;
    assign data_46 = data_43;
    assign data_48 = data_47;
    assign data_50 = data_49;
    assign data_52 = data_51;
    assign data_53 = data_51;
    assign data_54 = data_51;
    assign data_56 = data_55;
    assign data_57 = data_55;
    assign data_58 = data_55;
    assign data_60 = data_59;
    assign data_62 = data_61;
    assign data_64 = data_63;
    assign data_65 = data_63;
    assign data_66 = data_63;
    assign data_68 = data_67;
    assign data_69 = data_67;
    assign data_70 = data_67;
    assign data_72 = data_71;
    assign data_74 = data_73;
    assign data_76 = data_75;
    assign data_77 = data_75;
    assign data_78 = data_75;
    assign data_80 = data_79;
    assign data_81 = data_79;
    assign data_82 = data_79;
    assign data_84 = data_83;
    assign data_86 = data_85;
    assign data_88 = data_87;
    assign data_89 = data_87;
    assign data_90 = data_87;
    assign data_92 = data_91;
    assign data_93 = data_91;
    assign data_94 = data_91;

    /* output assignments */
    assign done_ = _1756;
    assign rd_q0 = _1755;
    assign rd_q1 = _1559;
    assign rd_q2 = _1363;
    assign rd_q3 = _1167;
    assign rd_q4 = _971;
    assign rd_q5 = _775;
    assign rd_q6 = _579;
    assign rd_q7 = _383;

endmodule
module multi_parallel_cores (
    rd_addr7,
    wr_addr7,
    wr_d_7_7,
    wr_d_7_6,
    wr_d_7_5,
    wr_d_7_4,
    wr_d_7_3,
    wr_d_7_2,
    wr_d_7_1,
    wr_d_7_0,
    rd_addr6,
    wr_addr6,
    wr_d_6_7,
    wr_d_6_6,
    wr_d_6_5,
    wr_d_6_4,
    wr_d_6_3,
    wr_d_6_2,
    wr_d_6_1,
    wr_d_6_0,
    rd_addr5,
    wr_addr5,
    wr_d_5_7,
    wr_d_5_6,
    wr_d_5_5,
    wr_d_5_4,
    wr_d_5_3,
    wr_d_5_2,
    wr_d_5_1,
    wr_d_5_0,
    rd_addr4,
    wr_addr4,
    wr_d_4_7,
    wr_d_4_6,
    wr_d_4_5,
    wr_d_4_4,
    wr_d_4_3,
    wr_d_4_2,
    wr_d_4_1,
    wr_d_4_0,
    rd_addr3,
    wr_addr3,
    wr_d_3_7,
    wr_d_3_6,
    wr_d_3_5,
    wr_d_3_4,
    wr_d_3_3,
    wr_d_3_2,
    wr_d_3_1,
    wr_d_3_0,
    rd_addr2,
    wr_addr2,
    wr_d_2_7,
    wr_d_2_6,
    wr_d_2_5,
    wr_d_2_4,
    wr_d_2_3,
    wr_d_2_2,
    wr_d_2_1,
    wr_d_2_0,
    rd_addr1,
    wr_addr1,
    wr_d_1_7,
    wr_d_1_6,
    wr_d_1_5,
    wr_d_1_4,
    wr_d_1_3,
    wr_d_1_2,
    wr_d_1_1,
    wr_d_1_0,
    rd_addr0,
    rd_en,
    wr_addr0,
    wr_en,
    wr_d_0_7,
    wr_d_0_6,
    wr_d_0_5,
    wr_d_0_4,
    wr_d_0_3,
    wr_d_0_2,
    wr_d_0_1,
    wr_d_0_0,
    flip,
    first_iter,
    first_4step_pass,
    start,
    clear,
    clock,
    done_,
    rd_d_0_0,
    rd_d_0_1,
    rd_d_0_2,
    rd_d_0_3,
    rd_d_0_4,
    rd_d_0_5,
    rd_d_0_6,
    rd_d_0_7,
    rd_d_1_0,
    rd_d_1_1,
    rd_d_1_2,
    rd_d_1_3,
    rd_d_1_4,
    rd_d_1_5,
    rd_d_1_6,
    rd_d_1_7,
    rd_d_2_0,
    rd_d_2_1,
    rd_d_2_2,
    rd_d_2_3,
    rd_d_2_4,
    rd_d_2_5,
    rd_d_2_6,
    rd_d_2_7,
    rd_d_3_0,
    rd_d_3_1,
    rd_d_3_2,
    rd_d_3_3,
    rd_d_3_4,
    rd_d_3_5,
    rd_d_3_6,
    rd_d_3_7,
    rd_d_4_0,
    rd_d_4_1,
    rd_d_4_2,
    rd_d_4_3,
    rd_d_4_4,
    rd_d_4_5,
    rd_d_4_6,
    rd_d_4_7,
    rd_d_5_0,
    rd_d_5_1,
    rd_d_5_2,
    rd_d_5_3,
    rd_d_5_4,
    rd_d_5_5,
    rd_d_5_6,
    rd_d_5_7,
    rd_d_6_0,
    rd_d_6_1,
    rd_d_6_2,
    rd_d_6_3,
    rd_d_6_4,
    rd_d_6_5,
    rd_d_6_6,
    rd_d_6_7,
    rd_d_7_0,
    rd_d_7_1,
    rd_d_7_2,
    rd_d_7_3,
    rd_d_7_4,
    rd_d_7_5,
    rd_d_7_6,
    rd_d_7_7
);

    input [11:0] rd_addr7;
    input [11:0] wr_addr7;
    input [63:0] wr_d_7_7;
    input [63:0] wr_d_7_6;
    input [63:0] wr_d_7_5;
    input [63:0] wr_d_7_4;
    input [63:0] wr_d_7_3;
    input [63:0] wr_d_7_2;
    input [63:0] wr_d_7_1;
    input [63:0] wr_d_7_0;
    input [11:0] rd_addr6;
    input [11:0] wr_addr6;
    input [63:0] wr_d_6_7;
    input [63:0] wr_d_6_6;
    input [63:0] wr_d_6_5;
    input [63:0] wr_d_6_4;
    input [63:0] wr_d_6_3;
    input [63:0] wr_d_6_2;
    input [63:0] wr_d_6_1;
    input [63:0] wr_d_6_0;
    input [11:0] rd_addr5;
    input [11:0] wr_addr5;
    input [63:0] wr_d_5_7;
    input [63:0] wr_d_5_6;
    input [63:0] wr_d_5_5;
    input [63:0] wr_d_5_4;
    input [63:0] wr_d_5_3;
    input [63:0] wr_d_5_2;
    input [63:0] wr_d_5_1;
    input [63:0] wr_d_5_0;
    input [11:0] rd_addr4;
    input [11:0] wr_addr4;
    input [63:0] wr_d_4_7;
    input [63:0] wr_d_4_6;
    input [63:0] wr_d_4_5;
    input [63:0] wr_d_4_4;
    input [63:0] wr_d_4_3;
    input [63:0] wr_d_4_2;
    input [63:0] wr_d_4_1;
    input [63:0] wr_d_4_0;
    input [11:0] rd_addr3;
    input [11:0] wr_addr3;
    input [63:0] wr_d_3_7;
    input [63:0] wr_d_3_6;
    input [63:0] wr_d_3_5;
    input [63:0] wr_d_3_4;
    input [63:0] wr_d_3_3;
    input [63:0] wr_d_3_2;
    input [63:0] wr_d_3_1;
    input [63:0] wr_d_3_0;
    input [11:0] rd_addr2;
    input [11:0] wr_addr2;
    input [63:0] wr_d_2_7;
    input [63:0] wr_d_2_6;
    input [63:0] wr_d_2_5;
    input [63:0] wr_d_2_4;
    input [63:0] wr_d_2_3;
    input [63:0] wr_d_2_2;
    input [63:0] wr_d_2_1;
    input [63:0] wr_d_2_0;
    input [11:0] rd_addr1;
    input [11:0] wr_addr1;
    input [63:0] wr_d_1_7;
    input [63:0] wr_d_1_6;
    input [63:0] wr_d_1_5;
    input [63:0] wr_d_1_4;
    input [63:0] wr_d_1_3;
    input [63:0] wr_d_1_2;
    input [63:0] wr_d_1_1;
    input [63:0] wr_d_1_0;
    input [11:0] rd_addr0;
    input [7:0] rd_en;
    input [11:0] wr_addr0;
    input [7:0] wr_en;
    input [63:0] wr_d_0_7;
    input [63:0] wr_d_0_6;
    input [63:0] wr_d_0_5;
    input [63:0] wr_d_0_4;
    input [63:0] wr_d_0_3;
    input [63:0] wr_d_0_2;
    input [63:0] wr_d_0_1;
    input [63:0] wr_d_0_0;
    input flip;
    input first_iter;
    input first_4step_pass;
    input start;
    input clear;
    input clock;
    output done_;
    output [63:0] rd_d_0_0;
    output [63:0] rd_d_0_1;
    output [63:0] rd_d_0_2;
    output [63:0] rd_d_0_3;
    output [63:0] rd_d_0_4;
    output [63:0] rd_d_0_5;
    output [63:0] rd_d_0_6;
    output [63:0] rd_d_0_7;
    output [63:0] rd_d_1_0;
    output [63:0] rd_d_1_1;
    output [63:0] rd_d_1_2;
    output [63:0] rd_d_1_3;
    output [63:0] rd_d_1_4;
    output [63:0] rd_d_1_5;
    output [63:0] rd_d_1_6;
    output [63:0] rd_d_1_7;
    output [63:0] rd_d_2_0;
    output [63:0] rd_d_2_1;
    output [63:0] rd_d_2_2;
    output [63:0] rd_d_2_3;
    output [63:0] rd_d_2_4;
    output [63:0] rd_d_2_5;
    output [63:0] rd_d_2_6;
    output [63:0] rd_d_2_7;
    output [63:0] rd_d_3_0;
    output [63:0] rd_d_3_1;
    output [63:0] rd_d_3_2;
    output [63:0] rd_d_3_3;
    output [63:0] rd_d_3_4;
    output [63:0] rd_d_3_5;
    output [63:0] rd_d_3_6;
    output [63:0] rd_d_3_7;
    output [63:0] rd_d_4_0;
    output [63:0] rd_d_4_1;
    output [63:0] rd_d_4_2;
    output [63:0] rd_d_4_3;
    output [63:0] rd_d_4_4;
    output [63:0] rd_d_4_5;
    output [63:0] rd_d_4_6;
    output [63:0] rd_d_4_7;
    output [63:0] rd_d_5_0;
    output [63:0] rd_d_5_1;
    output [63:0] rd_d_5_2;
    output [63:0] rd_d_5_3;
    output [63:0] rd_d_5_4;
    output [63:0] rd_d_5_5;
    output [63:0] rd_d_5_6;
    output [63:0] rd_d_5_7;
    output [63:0] rd_d_6_0;
    output [63:0] rd_d_6_1;
    output [63:0] rd_d_6_2;
    output [63:0] rd_d_6_3;
    output [63:0] rd_d_6_4;
    output [63:0] rd_d_6_5;
    output [63:0] rd_d_6_6;
    output [63:0] rd_d_6_7;
    output [63:0] rd_d_7_0;
    output [63:0] rd_d_7_1;
    output [63:0] rd_d_7_2;
    output [63:0] rd_d_7_3;
    output [63:0] rd_d_7_4;
    output [63:0] rd_d_7_5;
    output [63:0] rd_d_7_6;
    output [63:0] rd_d_7_7;

    /* signal declarations */
    wire [63:0] _252;
    wire [63:0] _253;
    wire [63:0] _254;
    wire [63:0] _255;
    wire [63:0] _256;
    wire [63:0] _257;
    wire [63:0] _258;
    wire [11:0] _9;
    wire _246;
    wire [1:0] _247;
    wire [3:0] _248;
    wire [7:0] _249;
    wire [11:0] _11;
    wire _242;
    wire [1:0] _243;
    wire [3:0] _244;
    wire [7:0] _245;
    wire [63:0] _13;
    wire [63:0] _15;
    wire [63:0] _17;
    wire [63:0] _19;
    wire [63:0] _21;
    wire [63:0] _23;
    wire [63:0] _25;
    wire [63:0] _27;
    wire [512:0] _251;
    wire [63:0] _259;
    wire [63:0] _270;
    wire [63:0] _271;
    wire [63:0] _272;
    wire [63:0] _273;
    wire [63:0] _274;
    wire [63:0] _275;
    wire [63:0] _276;
    wire [11:0] _37;
    wire _264;
    wire [1:0] _265;
    wire [3:0] _266;
    wire [7:0] _267;
    wire [11:0] _39;
    wire _260;
    wire [1:0] _261;
    wire [3:0] _262;
    wire [7:0] _263;
    wire [63:0] _41;
    wire [63:0] _43;
    wire [63:0] _45;
    wire [63:0] _47;
    wire [63:0] _49;
    wire [63:0] _51;
    wire [63:0] _53;
    wire [63:0] _55;
    wire [512:0] _269;
    wire [63:0] _277;
    wire [63:0] _288;
    wire [63:0] _289;
    wire [63:0] _290;
    wire [63:0] _291;
    wire [63:0] _292;
    wire [63:0] _293;
    wire [63:0] _294;
    wire [11:0] _65;
    wire _282;
    wire [1:0] _283;
    wire [3:0] _284;
    wire [7:0] _285;
    wire [11:0] _67;
    wire _278;
    wire [1:0] _279;
    wire [3:0] _280;
    wire [7:0] _281;
    wire [63:0] _69;
    wire [63:0] _71;
    wire [63:0] _73;
    wire [63:0] _75;
    wire [63:0] _77;
    wire [63:0] _79;
    wire [63:0] _81;
    wire [63:0] _83;
    wire [512:0] _287;
    wire [63:0] _295;
    wire [63:0] _306;
    wire [63:0] _307;
    wire [63:0] _308;
    wire [63:0] _309;
    wire [63:0] _310;
    wire [63:0] _311;
    wire [63:0] _312;
    wire [11:0] _93;
    wire _300;
    wire [1:0] _301;
    wire [3:0] _302;
    wire [7:0] _303;
    wire [11:0] _95;
    wire _296;
    wire [1:0] _297;
    wire [3:0] _298;
    wire [7:0] _299;
    wire [63:0] _97;
    wire [63:0] _99;
    wire [63:0] _101;
    wire [63:0] _103;
    wire [63:0] _105;
    wire [63:0] _107;
    wire [63:0] _109;
    wire [63:0] _111;
    wire [512:0] _305;
    wire [63:0] _313;
    wire [63:0] _324;
    wire [63:0] _325;
    wire [63:0] _326;
    wire [63:0] _327;
    wire [63:0] _328;
    wire [63:0] _329;
    wire [63:0] _330;
    wire [11:0] _121;
    wire _318;
    wire [1:0] _319;
    wire [3:0] _320;
    wire [7:0] _321;
    wire [11:0] _123;
    wire _314;
    wire [1:0] _315;
    wire [3:0] _316;
    wire [7:0] _317;
    wire [63:0] _125;
    wire [63:0] _127;
    wire [63:0] _129;
    wire [63:0] _131;
    wire [63:0] _133;
    wire [63:0] _135;
    wire [63:0] _137;
    wire [63:0] _139;
    wire [512:0] _323;
    wire [63:0] _331;
    wire [63:0] _342;
    wire [63:0] _343;
    wire [63:0] _344;
    wire [63:0] _345;
    wire [63:0] _346;
    wire [63:0] _347;
    wire [63:0] _348;
    wire [11:0] _149;
    wire _336;
    wire [1:0] _337;
    wire [3:0] _338;
    wire [7:0] _339;
    wire [11:0] _151;
    wire _332;
    wire [1:0] _333;
    wire [3:0] _334;
    wire [7:0] _335;
    wire [63:0] _153;
    wire [63:0] _155;
    wire [63:0] _157;
    wire [63:0] _159;
    wire [63:0] _161;
    wire [63:0] _163;
    wire [63:0] _165;
    wire [63:0] _167;
    wire [512:0] _341;
    wire [63:0] _349;
    wire [63:0] _360;
    wire [63:0] _361;
    wire [63:0] _362;
    wire [63:0] _363;
    wire [63:0] _364;
    wire [63:0] _365;
    wire [63:0] _366;
    wire [11:0] _177;
    wire _354;
    wire [1:0] _355;
    wire [3:0] _356;
    wire [7:0] _357;
    wire [11:0] _179;
    wire _350;
    wire [1:0] _351;
    wire [3:0] _352;
    wire [7:0] _353;
    wire [63:0] _181;
    wire [63:0] _183;
    wire [63:0] _185;
    wire [63:0] _187;
    wire [63:0] _189;
    wire [63:0] _191;
    wire [63:0] _193;
    wire [63:0] _195;
    wire [512:0] _359;
    wire [63:0] _367;
    wire [63:0] _378;
    wire [63:0] _379;
    wire [63:0] _380;
    wire [63:0] _381;
    wire [63:0] _382;
    wire [63:0] _383;
    wire [63:0] _384;
    wire [63:0] _385;
    wire [11:0] _206;
    wire [7:0] _208;
    wire _372;
    wire [1:0] _373;
    wire [3:0] _374;
    wire [7:0] _375;
    wire [11:0] _210;
    wire [7:0] _212;
    wire _368;
    wire [1:0] _369;
    wire [3:0] _370;
    wire [7:0] _371;
    wire [63:0] _214;
    wire [63:0] _216;
    wire [63:0] _218;
    wire [63:0] _220;
    wire [63:0] _222;
    wire [63:0] _224;
    wire [63:0] _226;
    wire [63:0] _228;
    wire _230;
    wire _232;
    wire _234;
    wire _236;
    wire _238;
    wire _240;
    wire [512:0] _377;
    wire _386;

    /* logic */
    assign _252 = _251[512:449];
    assign _253 = _251[448:385];
    assign _254 = _251[384:321];
    assign _255 = _251[320:257];
    assign _256 = _251[256:193];
    assign _257 = _251[192:129];
    assign _258 = _251[128:65];
    assign _9 = rd_addr7;
    assign _246 = _208[7:7];
    assign _247 = { _246, _246 };
    assign _248 = { _247, _247 };
    assign _249 = { _248, _248 };
    assign _11 = wr_addr7;
    assign _242 = _212[7:7];
    assign _243 = { _242, _242 };
    assign _244 = { _243, _243 };
    assign _245 = { _244, _244 };
    assign _13 = wr_d_7_7;
    assign _15 = wr_d_7_6;
    assign _17 = wr_d_7_5;
    assign _19 = wr_d_7_4;
    assign _21 = wr_d_7_3;
    assign _23 = wr_d_7_2;
    assign _25 = wr_d_7_1;
    assign _27 = wr_d_7_0;
    parallel_cores_6
        parallel_cores_6
        ( .clock(_240), .clear(_238), .start(_236), .first_4step_pass(_234), .first_iter(_232), .flip(_230), .wr_d0(_27), .wr_d1(_25), .wr_d2(_23), .wr_d3(_21), .wr_d4(_19), .wr_d5(_17), .wr_d6(_15), .wr_d7(_13), .wr_en(_245), .wr_addr(_11), .rd_en(_249), .rd_addr(_9), .rd_q7(_251[512:449]), .rd_q6(_251[448:385]), .rd_q5(_251[384:321]), .rd_q4(_251[320:257]), .rd_q3(_251[256:193]), .rd_q2(_251[192:129]), .rd_q1(_251[128:65]), .rd_q0(_251[64:1]), .done_(_251[0:0]) );
    assign _259 = _251[64:1];
    assign _270 = _269[512:449];
    assign _271 = _269[448:385];
    assign _272 = _269[384:321];
    assign _273 = _269[320:257];
    assign _274 = _269[256:193];
    assign _275 = _269[192:129];
    assign _276 = _269[128:65];
    assign _37 = rd_addr6;
    assign _264 = _208[6:6];
    assign _265 = { _264, _264 };
    assign _266 = { _265, _265 };
    assign _267 = { _266, _266 };
    assign _39 = wr_addr6;
    assign _260 = _212[6:6];
    assign _261 = { _260, _260 };
    assign _262 = { _261, _261 };
    assign _263 = { _262, _262 };
    assign _41 = wr_d_6_7;
    assign _43 = wr_d_6_6;
    assign _45 = wr_d_6_5;
    assign _47 = wr_d_6_4;
    assign _49 = wr_d_6_3;
    assign _51 = wr_d_6_2;
    assign _53 = wr_d_6_1;
    assign _55 = wr_d_6_0;
    parallel_cores_5
        parallel_cores_5
        ( .clock(_240), .clear(_238), .start(_236), .first_4step_pass(_234), .first_iter(_232), .flip(_230), .wr_d0(_55), .wr_d1(_53), .wr_d2(_51), .wr_d3(_49), .wr_d4(_47), .wr_d5(_45), .wr_d6(_43), .wr_d7(_41), .wr_en(_263), .wr_addr(_39), .rd_en(_267), .rd_addr(_37), .rd_q7(_269[512:449]), .rd_q6(_269[448:385]), .rd_q5(_269[384:321]), .rd_q4(_269[320:257]), .rd_q3(_269[256:193]), .rd_q2(_269[192:129]), .rd_q1(_269[128:65]), .rd_q0(_269[64:1]), .done_(_269[0:0]) );
    assign _277 = _269[64:1];
    assign _288 = _287[512:449];
    assign _289 = _287[448:385];
    assign _290 = _287[384:321];
    assign _291 = _287[320:257];
    assign _292 = _287[256:193];
    assign _293 = _287[192:129];
    assign _294 = _287[128:65];
    assign _65 = rd_addr5;
    assign _282 = _208[5:5];
    assign _283 = { _282, _282 };
    assign _284 = { _283, _283 };
    assign _285 = { _284, _284 };
    assign _67 = wr_addr5;
    assign _278 = _212[5:5];
    assign _279 = { _278, _278 };
    assign _280 = { _279, _279 };
    assign _281 = { _280, _280 };
    assign _69 = wr_d_5_7;
    assign _71 = wr_d_5_6;
    assign _73 = wr_d_5_5;
    assign _75 = wr_d_5_4;
    assign _77 = wr_d_5_3;
    assign _79 = wr_d_5_2;
    assign _81 = wr_d_5_1;
    assign _83 = wr_d_5_0;
    parallel_cores_4
        parallel_cores_4
        ( .clock(_240), .clear(_238), .start(_236), .first_4step_pass(_234), .first_iter(_232), .flip(_230), .wr_d0(_83), .wr_d1(_81), .wr_d2(_79), .wr_d3(_77), .wr_d4(_75), .wr_d5(_73), .wr_d6(_71), .wr_d7(_69), .wr_en(_281), .wr_addr(_67), .rd_en(_285), .rd_addr(_65), .rd_q7(_287[512:449]), .rd_q6(_287[448:385]), .rd_q5(_287[384:321]), .rd_q4(_287[320:257]), .rd_q3(_287[256:193]), .rd_q2(_287[192:129]), .rd_q1(_287[128:65]), .rd_q0(_287[64:1]), .done_(_287[0:0]) );
    assign _295 = _287[64:1];
    assign _306 = _305[512:449];
    assign _307 = _305[448:385];
    assign _308 = _305[384:321];
    assign _309 = _305[320:257];
    assign _310 = _305[256:193];
    assign _311 = _305[192:129];
    assign _312 = _305[128:65];
    assign _93 = rd_addr4;
    assign _300 = _208[4:4];
    assign _301 = { _300, _300 };
    assign _302 = { _301, _301 };
    assign _303 = { _302, _302 };
    assign _95 = wr_addr4;
    assign _296 = _212[4:4];
    assign _297 = { _296, _296 };
    assign _298 = { _297, _297 };
    assign _299 = { _298, _298 };
    assign _97 = wr_d_4_7;
    assign _99 = wr_d_4_6;
    assign _101 = wr_d_4_5;
    assign _103 = wr_d_4_4;
    assign _105 = wr_d_4_3;
    assign _107 = wr_d_4_2;
    assign _109 = wr_d_4_1;
    assign _111 = wr_d_4_0;
    parallel_cores_3
        parallel_cores_3
        ( .clock(_240), .clear(_238), .start(_236), .first_4step_pass(_234), .first_iter(_232), .flip(_230), .wr_d0(_111), .wr_d1(_109), .wr_d2(_107), .wr_d3(_105), .wr_d4(_103), .wr_d5(_101), .wr_d6(_99), .wr_d7(_97), .wr_en(_299), .wr_addr(_95), .rd_en(_303), .rd_addr(_93), .rd_q7(_305[512:449]), .rd_q6(_305[448:385]), .rd_q5(_305[384:321]), .rd_q4(_305[320:257]), .rd_q3(_305[256:193]), .rd_q2(_305[192:129]), .rd_q1(_305[128:65]), .rd_q0(_305[64:1]), .done_(_305[0:0]) );
    assign _313 = _305[64:1];
    assign _324 = _323[512:449];
    assign _325 = _323[448:385];
    assign _326 = _323[384:321];
    assign _327 = _323[320:257];
    assign _328 = _323[256:193];
    assign _329 = _323[192:129];
    assign _330 = _323[128:65];
    assign _121 = rd_addr3;
    assign _318 = _208[3:3];
    assign _319 = { _318, _318 };
    assign _320 = { _319, _319 };
    assign _321 = { _320, _320 };
    assign _123 = wr_addr3;
    assign _314 = _212[3:3];
    assign _315 = { _314, _314 };
    assign _316 = { _315, _315 };
    assign _317 = { _316, _316 };
    assign _125 = wr_d_3_7;
    assign _127 = wr_d_3_6;
    assign _129 = wr_d_3_5;
    assign _131 = wr_d_3_4;
    assign _133 = wr_d_3_3;
    assign _135 = wr_d_3_2;
    assign _137 = wr_d_3_1;
    assign _139 = wr_d_3_0;
    parallel_cores_2
        parallel_cores_2
        ( .clock(_240), .clear(_238), .start(_236), .first_4step_pass(_234), .first_iter(_232), .flip(_230), .wr_d0(_139), .wr_d1(_137), .wr_d2(_135), .wr_d3(_133), .wr_d4(_131), .wr_d5(_129), .wr_d6(_127), .wr_d7(_125), .wr_en(_317), .wr_addr(_123), .rd_en(_321), .rd_addr(_121), .rd_q7(_323[512:449]), .rd_q6(_323[448:385]), .rd_q5(_323[384:321]), .rd_q4(_323[320:257]), .rd_q3(_323[256:193]), .rd_q2(_323[192:129]), .rd_q1(_323[128:65]), .rd_q0(_323[64:1]), .done_(_323[0:0]) );
    assign _331 = _323[64:1];
    assign _342 = _341[512:449];
    assign _343 = _341[448:385];
    assign _344 = _341[384:321];
    assign _345 = _341[320:257];
    assign _346 = _341[256:193];
    assign _347 = _341[192:129];
    assign _348 = _341[128:65];
    assign _149 = rd_addr2;
    assign _336 = _208[2:2];
    assign _337 = { _336, _336 };
    assign _338 = { _337, _337 };
    assign _339 = { _338, _338 };
    assign _151 = wr_addr2;
    assign _332 = _212[2:2];
    assign _333 = { _332, _332 };
    assign _334 = { _333, _333 };
    assign _335 = { _334, _334 };
    assign _153 = wr_d_2_7;
    assign _155 = wr_d_2_6;
    assign _157 = wr_d_2_5;
    assign _159 = wr_d_2_4;
    assign _161 = wr_d_2_3;
    assign _163 = wr_d_2_2;
    assign _165 = wr_d_2_1;
    assign _167 = wr_d_2_0;
    parallel_cores_1
        parallel_cores_1
        ( .clock(_240), .clear(_238), .start(_236), .first_4step_pass(_234), .first_iter(_232), .flip(_230), .wr_d0(_167), .wr_d1(_165), .wr_d2(_163), .wr_d3(_161), .wr_d4(_159), .wr_d5(_157), .wr_d6(_155), .wr_d7(_153), .wr_en(_335), .wr_addr(_151), .rd_en(_339), .rd_addr(_149), .rd_q7(_341[512:449]), .rd_q6(_341[448:385]), .rd_q5(_341[384:321]), .rd_q4(_341[320:257]), .rd_q3(_341[256:193]), .rd_q2(_341[192:129]), .rd_q1(_341[128:65]), .rd_q0(_341[64:1]), .done_(_341[0:0]) );
    assign _349 = _341[64:1];
    assign _360 = _359[512:449];
    assign _361 = _359[448:385];
    assign _362 = _359[384:321];
    assign _363 = _359[320:257];
    assign _364 = _359[256:193];
    assign _365 = _359[192:129];
    assign _366 = _359[128:65];
    assign _177 = rd_addr1;
    assign _354 = _208[1:1];
    assign _355 = { _354, _354 };
    assign _356 = { _355, _355 };
    assign _357 = { _356, _356 };
    assign _179 = wr_addr1;
    assign _350 = _212[1:1];
    assign _351 = { _350, _350 };
    assign _352 = { _351, _351 };
    assign _353 = { _352, _352 };
    assign _181 = wr_d_1_7;
    assign _183 = wr_d_1_6;
    assign _185 = wr_d_1_5;
    assign _187 = wr_d_1_4;
    assign _189 = wr_d_1_3;
    assign _191 = wr_d_1_2;
    assign _193 = wr_d_1_1;
    assign _195 = wr_d_1_0;
    parallel_cores_0
        parallel_cores_0
        ( .clock(_240), .clear(_238), .start(_236), .first_4step_pass(_234), .first_iter(_232), .flip(_230), .wr_d0(_195), .wr_d1(_193), .wr_d2(_191), .wr_d3(_189), .wr_d4(_187), .wr_d5(_185), .wr_d6(_183), .wr_d7(_181), .wr_en(_353), .wr_addr(_179), .rd_en(_357), .rd_addr(_177), .rd_q7(_359[512:449]), .rd_q6(_359[448:385]), .rd_q5(_359[384:321]), .rd_q4(_359[320:257]), .rd_q3(_359[256:193]), .rd_q2(_359[192:129]), .rd_q1(_359[128:65]), .rd_q0(_359[64:1]), .done_(_359[0:0]) );
    assign _367 = _359[64:1];
    assign _378 = _377[512:449];
    assign _379 = _377[448:385];
    assign _380 = _377[384:321];
    assign _381 = _377[320:257];
    assign _382 = _377[256:193];
    assign _383 = _377[192:129];
    assign _384 = _377[128:65];
    assign _385 = _377[64:1];
    assign _206 = rd_addr0;
    assign _208 = rd_en;
    assign _372 = _208[0:0];
    assign _373 = { _372, _372 };
    assign _374 = { _373, _373 };
    assign _375 = { _374, _374 };
    assign _210 = wr_addr0;
    assign _212 = wr_en;
    assign _368 = _212[0:0];
    assign _369 = { _368, _368 };
    assign _370 = { _369, _369 };
    assign _371 = { _370, _370 };
    assign _214 = wr_d_0_7;
    assign _216 = wr_d_0_6;
    assign _218 = wr_d_0_5;
    assign _220 = wr_d_0_4;
    assign _222 = wr_d_0_3;
    assign _224 = wr_d_0_2;
    assign _226 = wr_d_0_1;
    assign _228 = wr_d_0_0;
    assign _230 = flip;
    assign _232 = first_iter;
    assign _234 = first_4step_pass;
    assign _236 = start;
    assign _238 = clear;
    assign _240 = clock;
    parallel_cores
        parallel_cores
        ( .clock(_240), .clear(_238), .start(_236), .first_4step_pass(_234), .first_iter(_232), .flip(_230), .wr_d0(_228), .wr_d1(_226), .wr_d2(_224), .wr_d3(_222), .wr_d4(_220), .wr_d5(_218), .wr_d6(_216), .wr_d7(_214), .wr_en(_371), .wr_addr(_210), .rd_en(_375), .rd_addr(_206), .rd_q7(_377[512:449]), .rd_q6(_377[448:385]), .rd_q5(_377[384:321]), .rd_q4(_377[320:257]), .rd_q3(_377[256:193]), .rd_q2(_377[192:129]), .rd_q1(_377[128:65]), .rd_q0(_377[64:1]), .done_(_377[0:0]) );
    assign _386 = _377[0:0];

    /* aliases */

    /* output assignments */
    assign done_ = _386;
    assign rd_d_0_0 = _385;
    assign rd_d_0_1 = _384;
    assign rd_d_0_2 = _383;
    assign rd_d_0_3 = _382;
    assign rd_d_0_4 = _381;
    assign rd_d_0_5 = _380;
    assign rd_d_0_6 = _379;
    assign rd_d_0_7 = _378;
    assign rd_d_1_0 = _367;
    assign rd_d_1_1 = _366;
    assign rd_d_1_2 = _365;
    assign rd_d_1_3 = _364;
    assign rd_d_1_4 = _363;
    assign rd_d_1_5 = _362;
    assign rd_d_1_6 = _361;
    assign rd_d_1_7 = _360;
    assign rd_d_2_0 = _349;
    assign rd_d_2_1 = _348;
    assign rd_d_2_2 = _347;
    assign rd_d_2_3 = _346;
    assign rd_d_2_4 = _345;
    assign rd_d_2_5 = _344;
    assign rd_d_2_6 = _343;
    assign rd_d_2_7 = _342;
    assign rd_d_3_0 = _331;
    assign rd_d_3_1 = _330;
    assign rd_d_3_2 = _329;
    assign rd_d_3_3 = _328;
    assign rd_d_3_4 = _327;
    assign rd_d_3_5 = _326;
    assign rd_d_3_6 = _325;
    assign rd_d_3_7 = _324;
    assign rd_d_4_0 = _313;
    assign rd_d_4_1 = _312;
    assign rd_d_4_2 = _311;
    assign rd_d_4_3 = _310;
    assign rd_d_4_4 = _309;
    assign rd_d_4_5 = _308;
    assign rd_d_4_6 = _307;
    assign rd_d_4_7 = _306;
    assign rd_d_5_0 = _295;
    assign rd_d_5_1 = _294;
    assign rd_d_5_2 = _293;
    assign rd_d_5_3 = _292;
    assign rd_d_5_4 = _291;
    assign rd_d_5_5 = _290;
    assign rd_d_5_6 = _289;
    assign rd_d_5_7 = _288;
    assign rd_d_6_0 = _277;
    assign rd_d_6_1 = _276;
    assign rd_d_6_2 = _275;
    assign rd_d_6_3 = _274;
    assign rd_d_6_4 = _273;
    assign rd_d_6_5 = _272;
    assign rd_d_6_6 = _271;
    assign rd_d_6_7 = _270;
    assign rd_d_7_0 = _259;
    assign rd_d_7_1 = _258;
    assign rd_d_7_2 = _257;
    assign rd_d_7_3 = _256;
    assign rd_d_7_4 = _255;
    assign rd_d_7_5 = _254;
    assign rd_d_7_6 = _253;
    assign rd_d_7_7 = _252;

endmodule
module kernel (
    data_in_tdata,
    data_in_tvalid,
    first_4step_pass,
    start,
    data_out_dest_tready,
    clear,
    clock,
    data_in_tkeep,
    data_in_tlast,
    data_in_tstrb,
    data_out_tvalid,
    data_out_tdata,
    data_out_tkeep,
    data_out_tstrb,
    data_out_tlast,
    data_in_dest_tready,
    done_
);

    input [511:0] data_in_tdata;
    input data_in_tvalid;
    input first_4step_pass;
    input start;
    input data_out_dest_tready;
    input clear;
    input clock;
    input [63:0] data_in_tkeep;
    input data_in_tlast;
    input [63:0] data_in_tstrb;
    output data_out_tvalid;
    output [511:0] data_out_tdata;
    output [63:0] data_out_tkeep;
    output [63:0] data_out_tstrb;
    output data_out_tlast;
    output data_in_dest_tready;
    output done_;

    /* signal declarations */
    wire _33;
    wire _34;
    wire gnd = 1'b0;
    wire [63:0] _36 = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    wire [63:0] _37 = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    wire [511:0] _377 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _376 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _374 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _373 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _370 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _369 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _367 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _366 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _364 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _363 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _361;
    wire [63:0] _360;
    wire [63:0] _359;
    wire [63:0] _358;
    wire [63:0] _357;
    wire [63:0] _356;
    wire [63:0] _355;
    wire [63:0] _354;
    wire [511:0] _362;
    (* keep="TRUE" *)
    reg [511:0] _365;
    (* keep="TRUE" *)
    reg [511:0] _368;
    (* keep="TRUE" *)
    reg [511:0] _371;
    wire [511:0] _352 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _351 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _349 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _348 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _346 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _345 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _343;
    wire [63:0] _342;
    wire [63:0] _341;
    wire [63:0] _340;
    wire [63:0] _339;
    wire [63:0] _338;
    wire [63:0] _337;
    wire [63:0] _336;
    wire [511:0] _344;
    (* keep="TRUE" *)
    reg [511:0] _347;
    (* keep="TRUE" *)
    reg [511:0] _350;
    (* keep="TRUE" *)
    reg [511:0] _353;
    wire [511:0] _334 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _333 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _331 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _330 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _328 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _327 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _325;
    wire [63:0] _324;
    wire [63:0] _323;
    wire [63:0] _322;
    wire [63:0] _321;
    wire [63:0] _320;
    wire [63:0] _319;
    wire [63:0] _318;
    wire [511:0] _326;
    (* keep="TRUE" *)
    reg [511:0] _329;
    (* keep="TRUE" *)
    reg [511:0] _332;
    (* keep="TRUE" *)
    reg [511:0] _335;
    wire [511:0] _316 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _315 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _313 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _312 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _310 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _309 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _307;
    wire [63:0] _306;
    wire [63:0] _305;
    wire [63:0] _304;
    wire [63:0] _303;
    wire [63:0] _302;
    wire [63:0] _301;
    wire [63:0] _300;
    wire [511:0] _308;
    (* keep="TRUE" *)
    reg [511:0] _311;
    (* keep="TRUE" *)
    reg [511:0] _314;
    (* keep="TRUE" *)
    reg [511:0] _317;
    wire [511:0] _298 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _297 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _295 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _294 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _292 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _291 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _289;
    wire [63:0] _288;
    wire [63:0] _287;
    wire [63:0] _286;
    wire [63:0] _285;
    wire [63:0] _284;
    wire [63:0] _283;
    wire [63:0] _282;
    wire [511:0] _290;
    (* keep="TRUE" *)
    reg [511:0] _293;
    (* keep="TRUE" *)
    reg [511:0] _296;
    (* keep="TRUE" *)
    reg [511:0] _299;
    wire [511:0] _280 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _279 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _277 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _276 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _274 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _273 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _271;
    wire [63:0] _270;
    wire [63:0] _269;
    wire [63:0] _268;
    wire [63:0] _267;
    wire [63:0] _266;
    wire [63:0] _265;
    wire [63:0] _264;
    wire [511:0] _272;
    (* keep="TRUE" *)
    reg [511:0] _275;
    (* keep="TRUE" *)
    reg [511:0] _278;
    (* keep="TRUE" *)
    reg [511:0] _281;
    wire [511:0] _262 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _261 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _259 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _258 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _256 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _255 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _253;
    wire [63:0] _252;
    wire [63:0] _251;
    wire [63:0] _250;
    wire [63:0] _249;
    wire [63:0] _248;
    wire [63:0] _247;
    wire [63:0] _246;
    wire [511:0] _254;
    (* keep="TRUE" *)
    reg [511:0] _257;
    (* keep="TRUE" *)
    reg [511:0] _260;
    (* keep="TRUE" *)
    reg [511:0] _263;
    wire [511:0] _244 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _243 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _241 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _240 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _238 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _237 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [63:0] _235;
    wire [63:0] _234;
    wire [63:0] _233;
    wire [63:0] _232;
    wire [63:0] _231;
    wire [63:0] _230;
    wire [63:0] _229;
    wire [63:0] _228;
    wire [511:0] _236;
    (* keep="TRUE" *)
    reg [511:0] _239;
    (* keep="TRUE" *)
    reg [511:0] _242;
    (* keep="TRUE" *)
    reg [511:0] _245;
    wire [2:0] _62 = 3'b000;
    wire [2:0] _61 = 3'b000;
    wire [2:0] _59 = 3'b000;
    wire [2:0] _58 = 3'b000;
    wire [2:0] _56 = 3'b000;
    wire [2:0] _55 = 3'b000;
    wire [2:0] _53 = 3'b000;
    wire [2:0] _52 = 3'b000;
    wire [2:0] _50 = 3'b000;
    wire [2:0] _49 = 3'b000;
    wire [2:0] _47 = 3'b000;
    wire [2:0] _46 = 3'b000;
    wire [7:0] _42 = 8'b00000000;
    wire _43;
    wire _44;
    wire [2:0] _40 = 3'b000;
    wire [2:0] _39 = 3'b000;
    wire [2:0] _38;
    reg [2:0] _45;
    reg [2:0] _48;
    reg [2:0] _51;
    reg [2:0] _54;
    reg [2:0] _57;
    reg [2:0] _60;
    reg [2:0] _63;
    reg [511:0] _372;
    reg [511:0] _375;
    reg [511:0] _378;
    wire [11:0] _224 = 12'b000000000000;
    wire [11:0] _223 = 12'b000000000000;
    wire [11:0] _221 = 12'b000000000000;
    wire [11:0] _220 = 12'b000000000000;
    wire [11:0] _218 = 12'b000000000000;
    wire [11:0] _217 = 12'b000000000000;
    (* keep="TRUE" *)
    reg [11:0] _219;
    (* keep="TRUE" *)
    reg [11:0] _222;
    (* keep="TRUE" *)
    reg [11:0] _225;
    wire [11:0] _215 = 12'b000000000000;
    wire [11:0] _214 = 12'b000000000000;
    wire [11:0] _212 = 12'b000000000000;
    wire [11:0] _211 = 12'b000000000000;
    wire [11:0] _209 = 12'b000000000000;
    wire [11:0] _208 = 12'b000000000000;
    (* keep="TRUE" *)
    reg [11:0] _210;
    (* keep="TRUE" *)
    reg [11:0] _213;
    (* keep="TRUE" *)
    reg [11:0] _216;
    wire [11:0] _206 = 12'b000000000000;
    wire [11:0] _205 = 12'b000000000000;
    wire [11:0] _203 = 12'b000000000000;
    wire [11:0] _202 = 12'b000000000000;
    wire [11:0] _200 = 12'b000000000000;
    wire [11:0] _199 = 12'b000000000000;
    (* keep="TRUE" *)
    reg [11:0] _201;
    (* keep="TRUE" *)
    reg [11:0] _204;
    (* keep="TRUE" *)
    reg [11:0] _207;
    wire [11:0] _197 = 12'b000000000000;
    wire [11:0] _196 = 12'b000000000000;
    wire [11:0] _194 = 12'b000000000000;
    wire [11:0] _193 = 12'b000000000000;
    wire [11:0] _191 = 12'b000000000000;
    wire [11:0] _190 = 12'b000000000000;
    (* keep="TRUE" *)
    reg [11:0] _192;
    (* keep="TRUE" *)
    reg [11:0] _195;
    (* keep="TRUE" *)
    reg [11:0] _198;
    wire [11:0] _188 = 12'b000000000000;
    wire [11:0] _187 = 12'b000000000000;
    wire [11:0] _185 = 12'b000000000000;
    wire [11:0] _184 = 12'b000000000000;
    wire [11:0] _182 = 12'b000000000000;
    wire [11:0] _181 = 12'b000000000000;
    (* keep="TRUE" *)
    reg [11:0] _183;
    (* keep="TRUE" *)
    reg [11:0] _186;
    (* keep="TRUE" *)
    reg [11:0] _189;
    wire [11:0] _179 = 12'b000000000000;
    wire [11:0] _178 = 12'b000000000000;
    wire [11:0] _176 = 12'b000000000000;
    wire [11:0] _175 = 12'b000000000000;
    wire [11:0] _173 = 12'b000000000000;
    wire [11:0] _172 = 12'b000000000000;
    (* keep="TRUE" *)
    reg [11:0] _174;
    (* keep="TRUE" *)
    reg [11:0] _177;
    (* keep="TRUE" *)
    reg [11:0] _180;
    wire [11:0] _170 = 12'b000000000000;
    wire [11:0] _169 = 12'b000000000000;
    wire [11:0] _167 = 12'b000000000000;
    wire [11:0] _166 = 12'b000000000000;
    wire [11:0] _164 = 12'b000000000000;
    wire [11:0] _163 = 12'b000000000000;
    (* keep="TRUE" *)
    reg [11:0] _165;
    (* keep="TRUE" *)
    reg [11:0] _168;
    (* keep="TRUE" *)
    reg [11:0] _171;
    wire [11:0] _161 = 12'b000000000000;
    wire [11:0] _160 = 12'b000000000000;
    wire [11:0] _158 = 12'b000000000000;
    wire [11:0] _157 = 12'b000000000000;
    wire [11:0] _155 = 12'b000000000000;
    wire [11:0] _154 = 12'b000000000000;
    wire [11:0] _153;
    (* keep="TRUE" *)
    reg [11:0] _156;
    (* keep="TRUE" *)
    reg [11:0] _159;
    (* keep="TRUE" *)
    reg [11:0] _162;
    wire [7:0] _151 = 8'b00000000;
    wire [7:0] _150 = 8'b00000000;
    wire [7:0] _148 = 8'b00000000;
    wire [7:0] _147 = 8'b00000000;
    wire [7:0] _145 = 8'b00000000;
    wire [7:0] _144 = 8'b00000000;
    wire [7:0] _41;
    (* keep="TRUE" *)
    reg [7:0] _146;
    (* keep="TRUE" *)
    reg [7:0] _149;
    (* keep="TRUE" *)
    reg [7:0] _152;
    wire [11:0] _142 = 12'b000000000000;
    wire [11:0] _141 = 12'b000000000000;
    wire [11:0] _139 = 12'b000000000000;
    wire [11:0] _138 = 12'b000000000000;
    (* keep="TRUE" *)
    reg [11:0] _140;
    (* keep="TRUE" *)
    reg [11:0] _143;
    wire [11:0] _136 = 12'b000000000000;
    wire [11:0] _135 = 12'b000000000000;
    wire [11:0] _133 = 12'b000000000000;
    wire [11:0] _132 = 12'b000000000000;
    (* keep="TRUE" *)
    reg [11:0] _134;
    (* keep="TRUE" *)
    reg [11:0] _137;
    wire [11:0] _130 = 12'b000000000000;
    wire [11:0] _129 = 12'b000000000000;
    wire [11:0] _127 = 12'b000000000000;
    wire [11:0] _126 = 12'b000000000000;
    (* keep="TRUE" *)
    reg [11:0] _128;
    (* keep="TRUE" *)
    reg [11:0] _131;
    wire [11:0] _124 = 12'b000000000000;
    wire [11:0] _123 = 12'b000000000000;
    wire [11:0] _121 = 12'b000000000000;
    wire [11:0] _120 = 12'b000000000000;
    (* keep="TRUE" *)
    reg [11:0] _122;
    (* keep="TRUE" *)
    reg [11:0] _125;
    wire [11:0] _118 = 12'b000000000000;
    wire [11:0] _117 = 12'b000000000000;
    wire [11:0] _115 = 12'b000000000000;
    wire [11:0] _114 = 12'b000000000000;
    (* keep="TRUE" *)
    reg [11:0] _116;
    (* keep="TRUE" *)
    reg [11:0] _119;
    wire [11:0] _112 = 12'b000000000000;
    wire [11:0] _111 = 12'b000000000000;
    wire [11:0] _109 = 12'b000000000000;
    wire [11:0] _108 = 12'b000000000000;
    (* keep="TRUE" *)
    reg [11:0] _110;
    (* keep="TRUE" *)
    reg [11:0] _113;
    wire [11:0] _106 = 12'b000000000000;
    wire [11:0] _105 = 12'b000000000000;
    wire [11:0] _103 = 12'b000000000000;
    wire [11:0] _102 = 12'b000000000000;
    (* keep="TRUE" *)
    reg [11:0] _104;
    (* keep="TRUE" *)
    reg [11:0] _107;
    wire [11:0] _100 = 12'b000000000000;
    wire [11:0] _99 = 12'b000000000000;
    wire [11:0] _97 = 12'b000000000000;
    wire [11:0] _96 = 12'b000000000000;
    wire [11:0] _95;
    (* keep="TRUE" *)
    reg [11:0] _98;
    (* keep="TRUE" *)
    reg [11:0] _101;
    wire [7:0] _93 = 8'b00000000;
    wire [7:0] _92 = 8'b00000000;
    wire [7:0] _90 = 8'b00000000;
    wire [7:0] _89 = 8'b00000000;
    wire [7:0] _88;
    (* keep="TRUE" *)
    reg [7:0] _91;
    (* keep="TRUE" *)
    reg [7:0] _94;
    wire [63:0] _87;
    wire [127:0] _85;
    wire [63:0] _86;
    wire [191:0] _83;
    wire [63:0] _84;
    wire [255:0] _81;
    wire [63:0] _82;
    wire [319:0] _79;
    wire [63:0] _80;
    wire [383:0] _77;
    wire [63:0] _78;
    wire [447:0] _75;
    wire [63:0] _76;
    wire [511:0] _72 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _71 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire vdd = 1'b1;
    wire [511:0] _68 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _67 = 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    wire [511:0] _8;
    reg [511:0] _70;
    reg [511:0] _73;
    wire [63:0] _74;
    wire _66;
    wire _65;
    wire _64;
    wire [4096:0] _227;
    wire _379;
    wire _9;
    wire _30;
    wire _380;
    wire _10;
    wire _12;
    wire _14;
    wire [21:0] _26;
    wire _27;
    wire _16;
    wire [5:0] _32;
    wire _381;
    wire _17;
    wire _19;
    wire _21;
    wire _23;
    wire [24:0] _29;
    wire _382;

    /* logic */
    assign _33 = _32[0:0];
    assign _34 = _26[1:1];
    assign _361 = _227[3648:3585];
    assign _360 = _227[3712:3649];
    assign _359 = _227[3776:3713];
    assign _358 = _227[3840:3777];
    assign _357 = _227[3904:3841];
    assign _356 = _227[3968:3905];
    assign _355 = _227[4032:3969];
    assign _354 = _227[4096:4033];
    assign _362 = { _354, _355, _356, _357, _358, _359, _360, _361 };
    always @(posedge _23) begin
        if (_44)
            _365 <= _362;
    end
    always @(posedge _23) begin
        if (_44)
            _368 <= _365;
    end
    always @(posedge _23) begin
        if (_44)
            _371 <= _368;
    end
    assign _343 = _227[3136:3073];
    assign _342 = _227[3200:3137];
    assign _341 = _227[3264:3201];
    assign _340 = _227[3328:3265];
    assign _339 = _227[3392:3329];
    assign _338 = _227[3456:3393];
    assign _337 = _227[3520:3457];
    assign _336 = _227[3584:3521];
    assign _344 = { _336, _337, _338, _339, _340, _341, _342, _343 };
    always @(posedge _23) begin
        if (_44)
            _347 <= _344;
    end
    always @(posedge _23) begin
        if (_44)
            _350 <= _347;
    end
    always @(posedge _23) begin
        if (_44)
            _353 <= _350;
    end
    assign _325 = _227[2624:2561];
    assign _324 = _227[2688:2625];
    assign _323 = _227[2752:2689];
    assign _322 = _227[2816:2753];
    assign _321 = _227[2880:2817];
    assign _320 = _227[2944:2881];
    assign _319 = _227[3008:2945];
    assign _318 = _227[3072:3009];
    assign _326 = { _318, _319, _320, _321, _322, _323, _324, _325 };
    always @(posedge _23) begin
        if (_44)
            _329 <= _326;
    end
    always @(posedge _23) begin
        if (_44)
            _332 <= _329;
    end
    always @(posedge _23) begin
        if (_44)
            _335 <= _332;
    end
    assign _307 = _227[2112:2049];
    assign _306 = _227[2176:2113];
    assign _305 = _227[2240:2177];
    assign _304 = _227[2304:2241];
    assign _303 = _227[2368:2305];
    assign _302 = _227[2432:2369];
    assign _301 = _227[2496:2433];
    assign _300 = _227[2560:2497];
    assign _308 = { _300, _301, _302, _303, _304, _305, _306, _307 };
    always @(posedge _23) begin
        if (_44)
            _311 <= _308;
    end
    always @(posedge _23) begin
        if (_44)
            _314 <= _311;
    end
    always @(posedge _23) begin
        if (_44)
            _317 <= _314;
    end
    assign _289 = _227[1600:1537];
    assign _288 = _227[1664:1601];
    assign _287 = _227[1728:1665];
    assign _286 = _227[1792:1729];
    assign _285 = _227[1856:1793];
    assign _284 = _227[1920:1857];
    assign _283 = _227[1984:1921];
    assign _282 = _227[2048:1985];
    assign _290 = { _282, _283, _284, _285, _286, _287, _288, _289 };
    always @(posedge _23) begin
        if (_44)
            _293 <= _290;
    end
    always @(posedge _23) begin
        if (_44)
            _296 <= _293;
    end
    always @(posedge _23) begin
        if (_44)
            _299 <= _296;
    end
    assign _271 = _227[1088:1025];
    assign _270 = _227[1152:1089];
    assign _269 = _227[1216:1153];
    assign _268 = _227[1280:1217];
    assign _267 = _227[1344:1281];
    assign _266 = _227[1408:1345];
    assign _265 = _227[1472:1409];
    assign _264 = _227[1536:1473];
    assign _272 = { _264, _265, _266, _267, _268, _269, _270, _271 };
    always @(posedge _23) begin
        if (_44)
            _275 <= _272;
    end
    always @(posedge _23) begin
        if (_44)
            _278 <= _275;
    end
    always @(posedge _23) begin
        if (_44)
            _281 <= _278;
    end
    assign _253 = _227[576:513];
    assign _252 = _227[640:577];
    assign _251 = _227[704:641];
    assign _250 = _227[768:705];
    assign _249 = _227[832:769];
    assign _248 = _227[896:833];
    assign _247 = _227[960:897];
    assign _246 = _227[1024:961];
    assign _254 = { _246, _247, _248, _249, _250, _251, _252, _253 };
    always @(posedge _23) begin
        if (_44)
            _257 <= _254;
    end
    always @(posedge _23) begin
        if (_44)
            _260 <= _257;
    end
    always @(posedge _23) begin
        if (_44)
            _263 <= _260;
    end
    assign _235 = _227[64:1];
    assign _234 = _227[128:65];
    assign _233 = _227[192:129];
    assign _232 = _227[256:193];
    assign _231 = _227[320:257];
    assign _230 = _227[384:321];
    assign _229 = _227[448:385];
    assign _228 = _227[512:449];
    assign _236 = { _228, _229, _230, _231, _232, _233, _234, _235 };
    always @(posedge _23) begin
        if (_44)
            _239 <= _236;
    end
    always @(posedge _23) begin
        if (_44)
            _242 <= _239;
    end
    always @(posedge _23) begin
        if (_44)
            _245 <= _242;
    end
    assign _43 = _41 == _42;
    assign _44 = ~ _43;
    assign _38 = _29[24:22];
    always @(posedge _23) begin
        if (_44)
            _45 <= _38;
    end
    always @(posedge _23) begin
        if (_44)
            _48 <= _45;
    end
    always @(posedge _23) begin
        if (_44)
            _51 <= _48;
    end
    always @(posedge _23) begin
        if (_44)
            _54 <= _51;
    end
    always @(posedge _23) begin
        if (_44)
            _57 <= _54;
    end
    always @(posedge _23) begin
        if (_44)
            _60 <= _57;
    end
    always @(posedge _23) begin
        if (_44)
            _63 <= _60;
    end
    always @* begin
        case (_63)
        0: _372 <= _245;
        1: _372 <= _263;
        2: _372 <= _281;
        3: _372 <= _299;
        4: _372 <= _317;
        5: _372 <= _335;
        6: _372 <= _353;
        default: _372 <= _371;
        endcase
    end
    always @(posedge _23) begin
        if (_44)
            _375 <= _372;
    end
    always @(posedge _23) begin
        if (_44)
            _378 <= _375;
    end
    always @(posedge _23) begin
        _219 <= _153;
    end
    always @(posedge _23) begin
        _222 <= _219;
    end
    always @(posedge _23) begin
        _225 <= _222;
    end
    always @(posedge _23) begin
        _210 <= _153;
    end
    always @(posedge _23) begin
        _213 <= _210;
    end
    always @(posedge _23) begin
        _216 <= _213;
    end
    always @(posedge _23) begin
        _201 <= _153;
    end
    always @(posedge _23) begin
        _204 <= _201;
    end
    always @(posedge _23) begin
        _207 <= _204;
    end
    always @(posedge _23) begin
        _192 <= _153;
    end
    always @(posedge _23) begin
        _195 <= _192;
    end
    always @(posedge _23) begin
        _198 <= _195;
    end
    always @(posedge _23) begin
        _183 <= _153;
    end
    always @(posedge _23) begin
        _186 <= _183;
    end
    always @(posedge _23) begin
        _189 <= _186;
    end
    always @(posedge _23) begin
        _174 <= _153;
    end
    always @(posedge _23) begin
        _177 <= _174;
    end
    always @(posedge _23) begin
        _180 <= _177;
    end
    always @(posedge _23) begin
        _165 <= _153;
    end
    always @(posedge _23) begin
        _168 <= _165;
    end
    always @(posedge _23) begin
        _171 <= _168;
    end
    assign _153 = _29[13:2];
    always @(posedge _23) begin
        _156 <= _153;
    end
    always @(posedge _23) begin
        _159 <= _156;
    end
    always @(posedge _23) begin
        _162 <= _159;
    end
    assign _41 = _29[21:14];
    always @(posedge _23) begin
        _146 <= _41;
    end
    always @(posedge _23) begin
        _149 <= _146;
    end
    always @(posedge _23) begin
        _152 <= _149;
    end
    always @(posedge _23) begin
        _140 <= _95;
    end
    always @(posedge _23) begin
        _143 <= _140;
    end
    always @(posedge _23) begin
        _134 <= _95;
    end
    always @(posedge _23) begin
        _137 <= _134;
    end
    always @(posedge _23) begin
        _128 <= _95;
    end
    always @(posedge _23) begin
        _131 <= _128;
    end
    always @(posedge _23) begin
        _122 <= _95;
    end
    always @(posedge _23) begin
        _125 <= _122;
    end
    always @(posedge _23) begin
        _116 <= _95;
    end
    always @(posedge _23) begin
        _119 <= _116;
    end
    always @(posedge _23) begin
        _110 <= _95;
    end
    always @(posedge _23) begin
        _113 <= _110;
    end
    always @(posedge _23) begin
        _104 <= _95;
    end
    always @(posedge _23) begin
        _107 <= _104;
    end
    assign _95 = _26[13:2];
    always @(posedge _23) begin
        _98 <= _95;
    end
    always @(posedge _23) begin
        _101 <= _98;
    end
    assign _88 = _26[21:14];
    always @(posedge _23) begin
        _91 <= _88;
    end
    always @(posedge _23) begin
        _94 <= _91;
    end
    assign _87 = _85[127:64];
    assign _85 = _83[191:64];
    assign _86 = _85[63:0];
    assign _83 = _81[255:64];
    assign _84 = _83[63:0];
    assign _81 = _79[319:64];
    assign _82 = _81[63:0];
    assign _79 = _77[383:64];
    assign _80 = _79[63:0];
    assign _77 = _75[447:64];
    assign _78 = _77[63:0];
    assign _75 = _73[511:64];
    assign _76 = _75[63:0];
    assign _8 = data_in_tdata;
    always @(posedge _23) begin
        _70 <= _8;
    end
    always @(posedge _23) begin
        _73 <= _70;
    end
    assign _74 = _73[63:0];
    assign _66 = _32[5:5];
    assign _65 = _32[4:4];
    assign _64 = _32[3:3];
    multi_parallel_cores
        multi_parallel_cores
        ( .clock(_23), .clear(_21), .start(_64), .first_4step_pass(_14), .first_iter(_65), .flip(_66), .wr_d_0_0(_74), .wr_d_0_1(_76), .wr_d_0_2(_78), .wr_d_0_3(_80), .wr_d_0_4(_82), .wr_d_0_5(_84), .wr_d_0_6(_86), .wr_d_0_7(_87), .wr_d_1_0(_74), .wr_d_1_1(_76), .wr_d_1_2(_78), .wr_d_1_3(_80), .wr_d_1_4(_82), .wr_d_1_5(_84), .wr_d_1_6(_86), .wr_d_1_7(_87), .wr_d_2_0(_74), .wr_d_2_1(_76), .wr_d_2_2(_78), .wr_d_2_3(_80), .wr_d_2_4(_82), .wr_d_2_5(_84), .wr_d_2_6(_86), .wr_d_2_7(_87), .wr_d_3_0(_74), .wr_d_3_1(_76), .wr_d_3_2(_78), .wr_d_3_3(_80), .wr_d_3_4(_82), .wr_d_3_5(_84), .wr_d_3_6(_86), .wr_d_3_7(_87), .wr_d_4_0(_74), .wr_d_4_1(_76), .wr_d_4_2(_78), .wr_d_4_3(_80), .wr_d_4_4(_82), .wr_d_4_5(_84), .wr_d_4_6(_86), .wr_d_4_7(_87), .wr_d_5_0(_74), .wr_d_5_1(_76), .wr_d_5_2(_78), .wr_d_5_3(_80), .wr_d_5_4(_82), .wr_d_5_5(_84), .wr_d_5_6(_86), .wr_d_5_7(_87), .wr_d_6_0(_74), .wr_d_6_1(_76), .wr_d_6_2(_78), .wr_d_6_3(_80), .wr_d_6_4(_82), .wr_d_6_5(_84), .wr_d_6_6(_86), .wr_d_6_7(_87), .wr_d_7_0(_74), .wr_d_7_1(_76), .wr_d_7_2(_78), .wr_d_7_3(_80), .wr_d_7_4(_82), .wr_d_7_5(_84), .wr_d_7_6(_86), .wr_d_7_7(_87), .wr_en(_94), .wr_addr0(_101), .wr_addr1(_107), .wr_addr2(_113), .wr_addr3(_119), .wr_addr4(_125), .wr_addr5(_131), .wr_addr6(_137), .wr_addr7(_143), .rd_en(_152), .rd_addr0(_162), .rd_addr1(_171), .rd_addr2(_180), .rd_addr3(_189), .rd_addr4(_198), .rd_addr5(_207), .rd_addr6(_216), .rd_addr7(_225), .rd_d_7_7(_227[4096:4033]), .rd_d_7_6(_227[4032:3969]), .rd_d_7_5(_227[3968:3905]), .rd_d_7_4(_227[3904:3841]), .rd_d_7_3(_227[3840:3777]), .rd_d_7_2(_227[3776:3713]), .rd_d_7_1(_227[3712:3649]), .rd_d_7_0(_227[3648:3585]), .rd_d_6_7(_227[3584:3521]), .rd_d_6_6(_227[3520:3457]), .rd_d_6_5(_227[3456:3393]), .rd_d_6_4(_227[3392:3329]), .rd_d_6_3(_227[3328:3265]), .rd_d_6_2(_227[3264:3201]), .rd_d_6_1(_227[3200:3137]), .rd_d_6_0(_227[3136:3073]), .rd_d_5_7(_227[3072:3009]), .rd_d_5_6(_227[3008:2945]), .rd_d_5_5(_227[2944:2881]), .rd_d_5_4(_227[2880:2817]), .rd_d_5_3(_227[2816:2753]), .rd_d_5_2(_227[2752:2689]), .rd_d_5_1(_227[2688:2625]), .rd_d_5_0(_227[2624:2561]), .rd_d_4_7(_227[2560:2497]), .rd_d_4_6(_227[2496:2433]), .rd_d_4_5(_227[2432:2369]), .rd_d_4_4(_227[2368:2305]), .rd_d_4_3(_227[2304:2241]), .rd_d_4_2(_227[2240:2177]), .rd_d_4_1(_227[2176:2113]), .rd_d_4_0(_227[2112:2049]), .rd_d_3_7(_227[2048:1985]), .rd_d_3_6(_227[1984:1921]), .rd_d_3_5(_227[1920:1857]), .rd_d_3_4(_227[1856:1793]), .rd_d_3_3(_227[1792:1729]), .rd_d_3_2(_227[1728:1665]), .rd_d_3_1(_227[1664:1601]), .rd_d_3_0(_227[1600:1537]), .rd_d_2_7(_227[1536:1473]), .rd_d_2_6(_227[1472:1409]), .rd_d_2_5(_227[1408:1345]), .rd_d_2_4(_227[1344:1281]), .rd_d_2_3(_227[1280:1217]), .rd_d_2_2(_227[1216:1153]), .rd_d_2_1(_227[1152:1089]), .rd_d_2_0(_227[1088:1025]), .rd_d_1_7(_227[1024:961]), .rd_d_1_6(_227[960:897]), .rd_d_1_5(_227[896:833]), .rd_d_1_4(_227[832:769]), .rd_d_1_3(_227[768:705]), .rd_d_1_2(_227[704:641]), .rd_d_1_1(_227[640:577]), .rd_d_1_0(_227[576:513]), .rd_d_0_7(_227[512:449]), .rd_d_0_6(_227[448:385]), .rd_d_0_5(_227[384:321]), .rd_d_0_4(_227[320:257]), .rd_d_0_3(_227[256:193]), .rd_d_0_2(_227[192:129]), .rd_d_0_1(_227[128:65]), .rd_d_0_0(_227[64:1]), .done_(_227[0:0]) );
    assign _379 = _227[0:0];
    assign _9 = _379;
    assign _30 = _29[0:0];
    assign _380 = _32[1:1];
    assign _10 = _380;
    assign _12 = data_in_tvalid;
    assign _14 = first_4step_pass;
    load_sm
        load_sm
        ( .clock(_23), .clear(_21), .first_4step_pass(_14), .tvalid(_12), .start(_10), .wr_en(_26[21:14]), .wr_addr(_26[13:2]), .tready(_26[1:1]), .done_(_26[0:0]) );
    assign _27 = _26[0:0];
    assign _16 = start;
    controller
        controller
        ( .clock(_23), .clear(_21), .start(_16), .input_done(_27), .output_done(_30), .cores_done(_9), .flip(_32[5:5]), .first_iter(_32[4:4]), .start_cores(_32[3:3]), .start_output(_32[2:2]), .start_input(_32[1:1]), .done_(_32[0:0]) );
    assign _381 = _32[2:2];
    assign _17 = _381;
    assign _19 = data_out_dest_tready;
    assign _21 = clear;
    assign _23 = clock;
    store_sm
        store_sm
        ( .clock(_23), .clear(_21), .tready(_19), .start(_17), .block(_29[24:22]), .rd_en(_29[21:14]), .rd_addr(_29[13:2]), .tvalid(_29[1:1]), .done_(_29[0:0]) );
    assign _382 = _29[1:1];

    /* aliases */

    /* output assignments */
    assign data_out_tvalid = _382;
    assign data_out_tdata = _378;
    assign data_out_tkeep = _37;
    assign data_out_tstrb = _36;
    assign data_out_tlast = gnd;
    assign data_in_dest_tready = _34;
    assign done_ = _33;

endmodule
module transposer_memories (
    write_enable,
    write_data,
    write_address,
    clock,
    read_address,
    read_data0,
    read_data1,
    read_data2,
    read_data3,
    read_data4,
    read_data5,
    read_data6,
    read_data7
);

    input [7:0] write_enable;
    input [511:0] write_data;
    input [3:0] write_address;
    input clock;
    input [3:0] read_address;
    (* RAM_STYLE="distributed" *)
    output [511:0] read_data0;
    (* RAM_STYLE="distributed" *)
    output [511:0] read_data1;
    (* RAM_STYLE="distributed" *)
    output [511:0] read_data2;
    (* RAM_STYLE="distributed" *)
    output [511:0] read_data3;
    (* RAM_STYLE="distributed" *)
    output [511:0] read_data4;
    (* RAM_STYLE="distributed" *)
    output [511:0] read_data5;
    (* RAM_STYLE="distributed" *)
    output [511:0] read_data6;
    (* RAM_STYLE="distributed" *)
    output [511:0] read_data7;

    /* signal declarations */
    wire _19;
    reg [511:0] _20[0:15];
    wire [511:0] _21;
    wire _22;
    reg [511:0] _23[0:15];
    wire [511:0] _24;
    wire _25;
    reg [511:0] _26[0:15];
    wire [511:0] _27;
    wire _28;
    reg [511:0] _29[0:15];
    wire [511:0] _30;
    wire _31;
    reg [511:0] _32[0:15];
    wire [511:0] _33;
    wire _34;
    reg [511:0] _35[0:15];
    wire [511:0] _36;
    wire _37;
    reg [511:0] _38[0:15];
    wire [511:0] _39;
    wire [7:0] _9;
    wire _40;
    wire [511:0] _11;
    wire [3:0] _13;
    wire _15;
    reg [511:0] _41[0:15];
    wire [3:0] _17;
    wire [511:0] _42;

    /* logic */
    assign _19 = _9[7:7];
    always @(posedge _15) begin
        if (_19)
            _20[_13] <= _11;
    end
    assign _21 = _20[_17];
    assign _22 = _9[6:6];
    always @(posedge _15) begin
        if (_22)
            _23[_13] <= _11;
    end
    assign _24 = _23[_17];
    assign _25 = _9[5:5];
    always @(posedge _15) begin
        if (_25)
            _26[_13] <= _11;
    end
    assign _27 = _26[_17];
    assign _28 = _9[4:4];
    always @(posedge _15) begin
        if (_28)
            _29[_13] <= _11;
    end
    assign _30 = _29[_17];
    assign _31 = _9[3:3];
    always @(posedge _15) begin
        if (_31)
            _32[_13] <= _11;
    end
    assign _33 = _32[_17];
    assign _34 = _9[2:2];
    always @(posedge _15) begin
        if (_34)
            _35[_13] <= _11;
    end
    assign _36 = _35[_17];
    assign _37 = _9[1:1];
    always @(posedge _15) begin
        if (_37)
            _38[_13] <= _11;
    end
    assign _39 = _38[_17];
    assign _9 = write_enable;
    assign _40 = _9[0:0];
    assign _11 = write_data;
    assign _13 = write_address;
    assign _15 = clock;
    always @(posedge _15) begin
        if (_40)
            _41[_13] <= _11;
    end
    assign _17 = read_address;
    assign _42 = _41[_17];

    /* aliases */

    /* output assignments */
    assign read_data0 = _42;
    assign read_data1 = _39;
    assign read_data2 = _36;
    assign read_data3 = _33;
    assign read_data4 = _30;
    assign read_data5 = _27;
    assign read_data6 = _24;
    assign read_data7 = _21;

endmodule
module transposer (
    in_tdata,
    in_tvalid,
    clear,
    clock,
    out_tready,
    in_tkeep,
    in_tlast,
    in_tstrb,
    out_tvalid,
    out_tdata,
    out_tkeep,
    out_tstrb,
    out_tlast,
    in_tready
);

    input [511:0] in_tdata;
    input in_tvalid;
    input clear;
    input clock;
    input out_tready;
    input [63:0] in_tkeep;
    input in_tlast;
    input [63:0] in_tstrb;
    output out_tvalid;
    output [511:0] out_tdata;
    output [63:0] out_tkeep;
    output [63:0] out_tstrb;
    output out_tlast;
    output in_tready;

    /* signal declarations */
    wire _48 = 1'b0;
    wire _47 = 1'b0;
    wire _72 = 1'b1;
    wire _73;
    wire _59 = 1'b0;
    wire _60;
    wire _61;
    wire _62;
    wire _46;
    wire _63;
    wire _44;
    wire _74;
    wire _1;
    reg _49;
    wire _2;
    wire gnd = 1'b0;
    wire _4;
    wire [63:0] _76 = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    wire [63:0] _6;
    wire [63:0] _77 = 64'b1111111111111111111111111111111111111111111111111111111111111111;
    wire [63:0] _8;
    wire [63:0] _225;
    wire [127:0] _223;
    wire [63:0] _224;
    wire [191:0] _221;
    wire [63:0] _222;
    wire [255:0] _219;
    wire [63:0] _220;
    wire [319:0] _217;
    wire [63:0] _218;
    wire [383:0] _215;
    wire [63:0] _216;
    wire [447:0] _213;
    wire [63:0] _214;
    wire [511:0] _211;
    wire [63:0] _212;
    reg [63:0] _226;
    wire [63:0] _209;
    wire [127:0] _207;
    wire [63:0] _208;
    wire [191:0] _205;
    wire [63:0] _206;
    wire [255:0] _203;
    wire [63:0] _204;
    wire [319:0] _201;
    wire [63:0] _202;
    wire [383:0] _199;
    wire [63:0] _200;
    wire [447:0] _197;
    wire [63:0] _198;
    wire [511:0] _195;
    wire [63:0] _196;
    reg [63:0] _210;
    wire [63:0] _193;
    wire [127:0] _191;
    wire [63:0] _192;
    wire [191:0] _189;
    wire [63:0] _190;
    wire [255:0] _187;
    wire [63:0] _188;
    wire [319:0] _185;
    wire [63:0] _186;
    wire [383:0] _183;
    wire [63:0] _184;
    wire [447:0] _181;
    wire [63:0] _182;
    wire [511:0] _179;
    wire [63:0] _180;
    reg [63:0] _194;
    wire [63:0] _177;
    wire [127:0] _175;
    wire [63:0] _176;
    wire [191:0] _173;
    wire [63:0] _174;
    wire [255:0] _171;
    wire [63:0] _172;
    wire [319:0] _169;
    wire [63:0] _170;
    wire [383:0] _167;
    wire [63:0] _168;
    wire [447:0] _165;
    wire [63:0] _166;
    wire [511:0] _163;
    wire [63:0] _164;
    reg [63:0] _178;
    wire [63:0] _161;
    wire [127:0] _159;
    wire [63:0] _160;
    wire [191:0] _157;
    wire [63:0] _158;
    wire [255:0] _155;
    wire [63:0] _156;
    wire [319:0] _153;
    wire [63:0] _154;
    wire [383:0] _151;
    wire [63:0] _152;
    wire [447:0] _149;
    wire [63:0] _150;
    wire [511:0] _147;
    wire [63:0] _148;
    reg [63:0] _162;
    wire [63:0] _145;
    wire [127:0] _143;
    wire [63:0] _144;
    wire [191:0] _141;
    wire [63:0] _142;
    wire [255:0] _139;
    wire [63:0] _140;
    wire [319:0] _137;
    wire [63:0] _138;
    wire [383:0] _135;
    wire [63:0] _136;
    wire [447:0] _133;
    wire [63:0] _134;
    wire [511:0] _131;
    wire [63:0] _132;
    reg [63:0] _146;
    wire [63:0] _129;
    wire [127:0] _127;
    wire [63:0] _128;
    wire [191:0] _125;
    wire [63:0] _126;
    wire [255:0] _123;
    wire [63:0] _124;
    wire [319:0] _121;
    wire [63:0] _122;
    wire [383:0] _119;
    wire [63:0] _120;
    wire [447:0] _117;
    wire [63:0] _118;
    wire [511:0] _115;
    wire [63:0] _116;
    reg [63:0] _130;
    wire [63:0] _113;
    wire [127:0] _111;
    wire [63:0] _112;
    wire [191:0] _109;
    wire [63:0] _110;
    wire [255:0] _107;
    wire [63:0] _108;
    wire [319:0] _105;
    wire [63:0] _106;
    wire [383:0] _103;
    wire [63:0] _104;
    wire [447:0] _101;
    wire [63:0] _102;
    wire [511:0] _11;
    wire [511:0] _12;
    wire _78;
    wire _79;
    wire [1:0] _80;
    wire [3:0] _81;
    wire [7:0] _82;
    wire [7:0] _83;
    wire [7:0] _13;
    wire _84;
    wire [3:0] _85;
    wire [3:0] _14;
    wire _89;
    wire [3:0] _93;
    wire [3:0] _15;
    wire [4095:0] _98;
    wire [511:0] _99;
    wire [63:0] _100;
    reg [63:0] _114;
    wire [511:0] _227;
    wire [511:0] _16;
    wire _314 = 1'b0;
    wire _313 = 1'b0;
    wire _321 = 1'b1;
    wire _322;
    wire _316 = 1'b0;
    wire _317;
    wire _318;
    wire _319;
    wire _312;
    wire _320;
    wire _265 = 1'b0;
    wire _264 = 1'b0;
    wire [1:0] _305 = 2'b10;
    wire [1:0] _306;
    wire _307;
    wire [1:0] _302 = 2'b01;
    wire [1:0] _65 = 2'b00;
    wire [1:0] _64 = 2'b00;
    wire [1:0] _258 = 2'b01;
    wire [1:0] _259;
    wire [1:0] _260;
    wire [1:0] _261;
    wire [1:0] _262;
    wire _40 = 1'b0;
    wire _39 = 1'b0;
    wire _255;
    wire [7:0] _56 = 8'b00000000;
    wire [7:0] _55 = 8'b00000000;
    wire [7:0] _239 = 8'b00000001;
    wire [7:0] _238 = 8'b00000000;
    wire [1:0] _68 = 2'b01;
    wire [1:0] _69;
    wire _70;
    wire [1:0] rd_pos;
    wire _67;
    wire _71;
    wire [7:0] _240;
    wire [7:0] _233 = 8'b00000000;
    wire _231 = 1'b0;
    wire [6:0] _230;
    wire [7:0] _232;
    wire [7:0] _234;
    wire [7:0] _235;
    wire [7:0] _236;
    wire _229;
    wire [7:0] _237;
    wire _228;
    wire [7:0] _241;
    wire [7:0] _19;
    reg [7:0] _57;
    wire _58;
    wire _251;
    wire [2:0] _53 = 3'b111;
    wire [2:0] _51 = 3'b000;
    wire [2:0] _50 = 3'b000;
    wire [2:0] _245 = 3'b000;
    wire [2:0] _243 = 3'b001;
    wire [2:0] _244;
    wire [2:0] _246;
    wire [2:0] _247;
    wire _242;
    wire [2:0] _248;
    wire [2:0] _20;
    reg [2:0] _52;
    wire _54;
    wire _252;
    wire _22;
    wire _253;
    wire _45 = 1'b1;
    wire _250;
    wire _254;
    wire _43 = 1'b0;
    wire _249;
    wire _256;
    wire _23;
    reg _42;
    wire _257;
    wire [1:0] _263;
    wire [1:0] _24;
    reg [1:0] _66;
    wire [1:0] wr_pos;
    wire [1:0] _303;
    wire [1:0] _87 = 2'b00;
    wire [1:0] _86 = 2'b00;
    wire [1:0] _273 = 2'b01;
    wire [1:0] _274;
    wire [1:0] _275;
    wire [1:0] _276;
    wire [1:0] _277;
    wire _268;
    wire [1:0] _278;
    wire [1:0] _26;
    reg [1:0] _88;
    wire _304;
    wire _308;
    wire _309;
    wire [2:0] _271 = 3'b111;
    wire [2:0] _91 = 3'b000;
    wire [2:0] _90 = 3'b000;
    wire [2:0] _289 = 3'b000;
    wire [2:0] _284 = 3'b000;
    wire [2:0] _282 = 3'b001;
    wire [2:0] _283;
    wire [2:0] _285;
    wire [2:0] _286;
    wire [2:0] _287;
    wire _281;
    wire [2:0] _288;
    wire _280;
    wire [2:0] _290;
    wire [2:0] _27;
    reg [2:0] _92;
    wire _272;
    wire _298;
    wire [2:0] _269 = 3'b111;
    wire vdd = 1'b1;
    wire [2:0] _95 = 3'b000;
    wire _29;
    wire [2:0] _94 = 3'b000;
    wire _31;
    wire [2:0] _292 = 3'b001;
    wire [2:0] _293;
    wire [2:0] _294;
    wire _291;
    wire [2:0] _295;
    wire [2:0] _32;
    reg [2:0] element_offset;
    wire _270;
    wire _299;
    wire _34;
    wire _300;
    wire _267 = 1'b1;
    wire _297;
    wire _301;
    wire _279 = 1'b0;
    wire _296;
    wire _310;
    wire _35;
    reg _266;
    wire _311;
    wire _323;
    wire _36;
    reg _315;
    wire _37;

    /* logic */
    assign _73 = _71 ? _72 : _49;
    assign _60 = _58 ? _59 : _49;
    assign _61 = _54 ? _60 : _49;
    assign _62 = _22 ? _61 : _49;
    assign _46 = _42 == _45;
    assign _63 = _46 ? _62 : _49;
    assign _44 = _42 == _43;
    assign _74 = _44 ? _73 : _63;
    assign _1 = _74;
    always @(posedge _31) begin
        if (_29)
            _49 <= _48;
        else
            _49 <= _1;
    end
    assign _2 = _49;
    assign _4 = gnd;
    assign _6 = _76;
    assign _8 = _77;
    assign _225 = _223[127:64];
    assign _223 = _221[191:64];
    assign _224 = _223[63:0];
    assign _221 = _219[255:64];
    assign _222 = _221[63:0];
    assign _219 = _217[319:64];
    assign _220 = _219[63:0];
    assign _217 = _215[383:64];
    assign _218 = _217[63:0];
    assign _215 = _213[447:64];
    assign _216 = _215[63:0];
    assign _213 = _211[511:64];
    assign _214 = _213[63:0];
    assign _211 = _98[511:0];
    assign _212 = _211[63:0];
    always @* begin
        case (element_offset)
        0: _226 <= _212;
        1: _226 <= _214;
        2: _226 <= _216;
        3: _226 <= _218;
        4: _226 <= _220;
        5: _226 <= _222;
        6: _226 <= _224;
        default: _226 <= _225;
        endcase
    end
    assign _209 = _207[127:64];
    assign _207 = _205[191:64];
    assign _208 = _207[63:0];
    assign _205 = _203[255:64];
    assign _206 = _205[63:0];
    assign _203 = _201[319:64];
    assign _204 = _203[63:0];
    assign _201 = _199[383:64];
    assign _202 = _201[63:0];
    assign _199 = _197[447:64];
    assign _200 = _199[63:0];
    assign _197 = _195[511:64];
    assign _198 = _197[63:0];
    assign _195 = _98[1023:512];
    assign _196 = _195[63:0];
    always @* begin
        case (element_offset)
        0: _210 <= _196;
        1: _210 <= _198;
        2: _210 <= _200;
        3: _210 <= _202;
        4: _210 <= _204;
        5: _210 <= _206;
        6: _210 <= _208;
        default: _210 <= _209;
        endcase
    end
    assign _193 = _191[127:64];
    assign _191 = _189[191:64];
    assign _192 = _191[63:0];
    assign _189 = _187[255:64];
    assign _190 = _189[63:0];
    assign _187 = _185[319:64];
    assign _188 = _187[63:0];
    assign _185 = _183[383:64];
    assign _186 = _185[63:0];
    assign _183 = _181[447:64];
    assign _184 = _183[63:0];
    assign _181 = _179[511:64];
    assign _182 = _181[63:0];
    assign _179 = _98[1535:1024];
    assign _180 = _179[63:0];
    always @* begin
        case (element_offset)
        0: _194 <= _180;
        1: _194 <= _182;
        2: _194 <= _184;
        3: _194 <= _186;
        4: _194 <= _188;
        5: _194 <= _190;
        6: _194 <= _192;
        default: _194 <= _193;
        endcase
    end
    assign _177 = _175[127:64];
    assign _175 = _173[191:64];
    assign _176 = _175[63:0];
    assign _173 = _171[255:64];
    assign _174 = _173[63:0];
    assign _171 = _169[319:64];
    assign _172 = _171[63:0];
    assign _169 = _167[383:64];
    assign _170 = _169[63:0];
    assign _167 = _165[447:64];
    assign _168 = _167[63:0];
    assign _165 = _163[511:64];
    assign _166 = _165[63:0];
    assign _163 = _98[2047:1536];
    assign _164 = _163[63:0];
    always @* begin
        case (element_offset)
        0: _178 <= _164;
        1: _178 <= _166;
        2: _178 <= _168;
        3: _178 <= _170;
        4: _178 <= _172;
        5: _178 <= _174;
        6: _178 <= _176;
        default: _178 <= _177;
        endcase
    end
    assign _161 = _159[127:64];
    assign _159 = _157[191:64];
    assign _160 = _159[63:0];
    assign _157 = _155[255:64];
    assign _158 = _157[63:0];
    assign _155 = _153[319:64];
    assign _156 = _155[63:0];
    assign _153 = _151[383:64];
    assign _154 = _153[63:0];
    assign _151 = _149[447:64];
    assign _152 = _151[63:0];
    assign _149 = _147[511:64];
    assign _150 = _149[63:0];
    assign _147 = _98[2559:2048];
    assign _148 = _147[63:0];
    always @* begin
        case (element_offset)
        0: _162 <= _148;
        1: _162 <= _150;
        2: _162 <= _152;
        3: _162 <= _154;
        4: _162 <= _156;
        5: _162 <= _158;
        6: _162 <= _160;
        default: _162 <= _161;
        endcase
    end
    assign _145 = _143[127:64];
    assign _143 = _141[191:64];
    assign _144 = _143[63:0];
    assign _141 = _139[255:64];
    assign _142 = _141[63:0];
    assign _139 = _137[319:64];
    assign _140 = _139[63:0];
    assign _137 = _135[383:64];
    assign _138 = _137[63:0];
    assign _135 = _133[447:64];
    assign _136 = _135[63:0];
    assign _133 = _131[511:64];
    assign _134 = _133[63:0];
    assign _131 = _98[3071:2560];
    assign _132 = _131[63:0];
    always @* begin
        case (element_offset)
        0: _146 <= _132;
        1: _146 <= _134;
        2: _146 <= _136;
        3: _146 <= _138;
        4: _146 <= _140;
        5: _146 <= _142;
        6: _146 <= _144;
        default: _146 <= _145;
        endcase
    end
    assign _129 = _127[127:64];
    assign _127 = _125[191:64];
    assign _128 = _127[63:0];
    assign _125 = _123[255:64];
    assign _126 = _125[63:0];
    assign _123 = _121[319:64];
    assign _124 = _123[63:0];
    assign _121 = _119[383:64];
    assign _122 = _121[63:0];
    assign _119 = _117[447:64];
    assign _120 = _119[63:0];
    assign _117 = _115[511:64];
    assign _118 = _117[63:0];
    assign _115 = _98[3583:3072];
    assign _116 = _115[63:0];
    always @* begin
        case (element_offset)
        0: _130 <= _116;
        1: _130 <= _118;
        2: _130 <= _120;
        3: _130 <= _122;
        4: _130 <= _124;
        5: _130 <= _126;
        6: _130 <= _128;
        default: _130 <= _129;
        endcase
    end
    assign _113 = _111[127:64];
    assign _111 = _109[191:64];
    assign _112 = _111[63:0];
    assign _109 = _107[255:64];
    assign _110 = _109[63:0];
    assign _107 = _105[319:64];
    assign _108 = _107[63:0];
    assign _105 = _103[383:64];
    assign _106 = _105[63:0];
    assign _103 = _101[447:64];
    assign _104 = _103[63:0];
    assign _101 = _99[511:64];
    assign _102 = _101[63:0];
    assign _11 = in_tdata;
    assign _12 = _11;
    assign _78 = _45 == _42;
    assign _79 = _78 & _22;
    assign _80 = { _79, _79 };
    assign _81 = { _80, _80 };
    assign _82 = { _81, _81 };
    assign _83 = _57 & _82;
    assign _13 = _83;
    assign _84 = _66[0:0];
    assign _85 = { _84, _52 };
    assign _14 = _85;
    assign _89 = _88[0:0];
    assign _93 = { _89, _92 };
    assign _15 = _93;
    transposer_memories
        transposer_memories
        ( .clock(_31), .read_address(_15), .write_address(_14), .write_enable(_13), .write_data(_12), .read_data7(_98[4095:3584]), .read_data6(_98[3583:3072]), .read_data5(_98[3071:2560]), .read_data4(_98[2559:2048]), .read_data3(_98[2047:1536]), .read_data2(_98[1535:1024]), .read_data1(_98[1023:512]), .read_data0(_98[511:0]) );
    assign _99 = _98[4095:3584];
    assign _100 = _99[63:0];
    always @* begin
        case (element_offset)
        0: _114 <= _100;
        1: _114 <= _102;
        2: _114 <= _104;
        3: _114 <= _106;
        4: _114 <= _108;
        5: _114 <= _110;
        6: _114 <= _112;
        default: _114 <= _113;
        endcase
    end
    assign _227 = { _114, _130, _146, _162, _178, _194, _210, _226 };
    assign _16 = _227;
    assign _322 = _308 ? _321 : _315;
    assign _317 = _272 ? _316 : _315;
    assign _318 = _270 ? _317 : _315;
    assign _319 = _34 ? _318 : _315;
    assign _312 = _266 == _267;
    assign _320 = _312 ? _319 : _315;
    assign _306 = wr_pos - _305;
    assign _307 = _88 == _306;
    assign _259 = _66 + _258;
    assign _260 = _58 ? _259 : _66;
    assign _261 = _54 ? _260 : _66;
    assign _262 = _22 ? _261 : _66;
    assign _255 = _71 ? _45 : _42;
    assign _69 = _66 - _68;
    assign _70 = rd_pos == _69;
    assign rd_pos = _88;
    assign _67 = rd_pos == _66;
    assign _71 = _67 | _70;
    assign _240 = _71 ? _239 : _238;
    assign _230 = _57[6:0];
    assign _232 = { _230, _231 };
    assign _234 = _58 ? _233 : _232;
    assign _235 = _54 ? _234 : _57;
    assign _236 = _22 ? _235 : _57;
    assign _229 = _42 == _45;
    assign _237 = _229 ? _236 : _57;
    assign _228 = _42 == _43;
    assign _241 = _228 ? _240 : _237;
    assign _19 = _241;
    always @(posedge _31) begin
        if (_29)
            _57 <= _56;
        else
            _57 <= _19;
    end
    assign _58 = _57[7:7];
    assign _251 = _58 ? _43 : _42;
    assign _244 = _52 + _243;
    assign _246 = _54 ? _245 : _244;
    assign _247 = _22 ? _246 : _52;
    assign _242 = _42 == _45;
    assign _248 = _242 ? _247 : _52;
    assign _20 = _248;
    always @(posedge _31) begin
        if (_29)
            _52 <= _51;
        else
            _52 <= _20;
    end
    assign _54 = _52 == _53;
    assign _252 = _54 ? _251 : _42;
    assign _22 = in_tvalid;
    assign _253 = _22 ? _252 : _42;
    assign _250 = _42 == _45;
    assign _254 = _250 ? _253 : _42;
    assign _249 = _42 == _43;
    assign _256 = _249 ? _255 : _254;
    assign _23 = _256;
    always @(posedge _31) begin
        if (_29)
            _42 <= _40;
        else
            _42 <= _23;
    end
    assign _257 = _42 == _45;
    assign _263 = _257 ? _262 : _66;
    assign _24 = _263;
    always @(posedge _31) begin
        if (_29)
            _66 <= _65;
        else
            _66 <= _24;
    end
    assign wr_pos = _66;
    assign _303 = wr_pos - _302;
    assign _274 = _88 + _273;
    assign _275 = _272 ? _274 : _88;
    assign _276 = _270 ? _275 : _88;
    assign _277 = _34 ? _276 : _88;
    assign _268 = _266 == _267;
    assign _278 = _268 ? _277 : _88;
    assign _26 = _278;
    always @(posedge _31) begin
        if (_29)
            _88 <= _87;
        else
            _88 <= _26;
    end
    assign _304 = _88 == _303;
    assign _308 = _304 | _307;
    assign _309 = _308 ? _267 : _266;
    assign _283 = _92 + _282;
    assign _285 = _272 ? _284 : _283;
    assign _286 = _270 ? _285 : _92;
    assign _287 = _34 ? _286 : _92;
    assign _281 = _266 == _267;
    assign _288 = _281 ? _287 : _92;
    assign _280 = _266 == _279;
    assign _290 = _280 ? _289 : _288;
    assign _27 = _290;
    always @(posedge _31) begin
        if (_29)
            _92 <= _91;
        else
            _92 <= _27;
    end
    assign _272 = _92 == _271;
    assign _298 = _272 ? _279 : _266;
    assign _29 = clear;
    assign _31 = clock;
    assign _293 = element_offset + _292;
    assign _294 = _34 ? _293 : element_offset;
    assign _291 = _266 == _267;
    assign _295 = _291 ? _294 : element_offset;
    assign _32 = _295;
    always @(posedge _31) begin
        if (_29)
            element_offset <= _95;
        else
            element_offset <= _32;
    end
    assign _270 = element_offset == _269;
    assign _299 = _270 ? _298 : _266;
    assign _34 = out_tready;
    assign _300 = _34 ? _299 : _266;
    assign _297 = _266 == _267;
    assign _301 = _297 ? _300 : _266;
    assign _296 = _266 == _279;
    assign _310 = _296 ? _309 : _301;
    assign _35 = _310;
    always @(posedge _31) begin
        if (_29)
            _266 <= _265;
        else
            _266 <= _35;
    end
    assign _311 = _266 == _279;
    assign _323 = _311 ? _322 : _320;
    assign _36 = _323;
    always @(posedge _31) begin
        if (_29)
            _315 <= _314;
        else
            _315 <= _36;
    end
    assign _37 = _315;

    /* aliases */

    /* output assignments */
    assign out_tvalid = _37;
    assign out_tdata = _16;
    assign out_tkeep = _8;
    assign out_tstrb = _6;
    assign out_tlast = _4;
    assign in_tready = _2;

endmodule
module krnl_ntt (
    compute_to_controller_tready,
    controller_to_compute_phase_1_tlast,
    controller_to_compute_phase_1_tstrb,
    controller_to_compute_phase_1_tkeep,
    controller_to_compute_phase_1_tdata,
    controller_to_compute_phase_2_tlast,
    controller_to_compute_phase_2_tstrb,
    controller_to_compute_phase_2_tkeep,
    controller_to_compute_phase_2_tdata,
    controller_to_compute_phase_2_tvalid,
    controller_to_compute_phase_1_tvalid,
    ap_rst_n,
    ap_clk,
    compute_to_controller_tvalid,
    compute_to_controller_tdata,
    compute_to_controller_tkeep,
    compute_to_controller_tstrb,
    compute_to_controller_tlast,
    controller_to_compute_phase_1_tready,
    controller_to_compute_phase_2_tready
);

    input compute_to_controller_tready;
    input controller_to_compute_phase_1_tlast;
    input [63:0] controller_to_compute_phase_1_tstrb;
    input [63:0] controller_to_compute_phase_1_tkeep;
    input [511:0] controller_to_compute_phase_1_tdata;
    input controller_to_compute_phase_2_tlast;
    input [63:0] controller_to_compute_phase_2_tstrb;
    input [63:0] controller_to_compute_phase_2_tkeep;
    input [511:0] controller_to_compute_phase_2_tdata;
    input controller_to_compute_phase_2_tvalid;
    input controller_to_compute_phase_1_tvalid;
    input ap_rst_n;
    input ap_clk;
    output compute_to_controller_tvalid;
    output [511:0] compute_to_controller_tdata;
    output [63:0] compute_to_controller_tkeep;
    output [63:0] compute_to_controller_tstrb;
    output compute_to_controller_tlast;
    output controller_to_compute_phase_1_tready;
    output controller_to_compute_phase_2_tready;

    /* signal declarations */
    wire _41;
    wire _57;
    wire [63:0] _58;
    wire [63:0] _59;
    wire [511:0] _60;
    wire _8;
    wire _10;
    wire _53;
    wire _54;
    wire [63:0] _12;
    wire [63:0] _51;
    wire [63:0] _52;
    wire [63:0] _14;
    wire [63:0] _49;
    wire [63:0] _50;
    wire [511:0] _16;
    wire [511:0] _47;
    wire [511:0] _48;
    wire _61;
    wire _17;
    wire _18;
    wire _20;
    wire [63:0] _22;
    wire [63:0] _24;
    wire [511:0] _26;
    wire [642:0] _40;
    wire _45;
    wire _46;
    wire _43 = 1'b0;
    wire _42 = 1'b0;
    wire _62;
    wire _27;
    reg _4STEP;
    wire _29;
    wire _31;
    wire _64;
    wire _63;
    wire _65;
    wire _32;
    wire _34;
    wire _38;
    wire _36;
    wire [643:0] _56;
    wire _66;

    /* logic */
    assign _41 = _40[642:642];
    assign _57 = _56[641:641];
    assign _58 = _56[640:577];
    assign _59 = _56[576:513];
    assign _60 = _56[512:1];
    assign _8 = compute_to_controller_tready;
    assign _10 = controller_to_compute_phase_1_tlast;
    assign _53 = _40[641:641];
    assign _54 = _31 ? _10 : _53;
    assign _12 = controller_to_compute_phase_1_tstrb;
    assign _51 = _40[640:577];
    assign _52 = _31 ? _12 : _51;
    assign _14 = controller_to_compute_phase_1_tkeep;
    assign _49 = _40[576:513];
    assign _50 = _31 ? _14 : _49;
    assign _16 = controller_to_compute_phase_1_tdata;
    assign _47 = _40[512:1];
    assign _48 = _31 ? _16 : _47;
    assign _61 = _56[642:642];
    assign _17 = _61;
    assign _18 = _17;
    assign _20 = controller_to_compute_phase_2_tlast;
    assign _22 = controller_to_compute_phase_2_tstrb;
    assign _24 = controller_to_compute_phase_2_tkeep;
    assign _26 = controller_to_compute_phase_2_tdata;
    transposer
        transposer
        ( .clock(_36), .clear(_38), .in_tvalid(_29), .in_tdata(_26), .in_tkeep(_24), .in_tstrb(_22), .in_tlast(_20), .out_tready(_18), .in_tready(_40[642:642]), .out_tlast(_40[641:641]), .out_tstrb(_40[640:577]), .out_tkeep(_40[576:513]), .out_tdata(_40[512:1]), .out_tvalid(_40[0:0]) );
    assign _45 = _40[0:0];
    assign _46 = _31 ? _31 : _45;
    assign _62 = ~ _4STEP;
    assign _27 = _62;
    always @(posedge _36) begin
        if (_38)
            _4STEP <= _43;
        else
            if (_32)
                _4STEP <= _27;
    end
    assign _29 = controller_to_compute_phase_2_tvalid;
    assign _31 = controller_to_compute_phase_1_tvalid;
    assign _64 = _31 | _29;
    assign _63 = _56[643:643];
    assign _65 = _63 & _64;
    assign _32 = _65;
    assign _34 = ap_rst_n;
    assign _38 = ~ _34;
    assign _36 = ap_clk;
    kernel
        kernel
        ( .clock(_36), .clear(_38), .start(_32), .first_4step_pass(_4STEP), .data_in_tvalid(_46), .data_in_tdata(_48), .data_in_tkeep(_50), .data_in_tstrb(_52), .data_in_tlast(_54), .data_out_dest_tready(_8), .done_(_56[643:643]), .data_in_dest_tready(_56[642:642]), .data_out_tlast(_56[641:641]), .data_out_tstrb(_56[640:577]), .data_out_tkeep(_56[576:513]), .data_out_tdata(_56[512:1]), .data_out_tvalid(_56[0:0]) );
    assign _66 = _56[0:0];

    /* aliases */

    /* output assignments */
    assign compute_to_controller_tvalid = _66;
    assign compute_to_controller_tdata = _60;
    assign compute_to_controller_tkeep = _59;
    assign compute_to_controller_tstrb = _58;
    assign compute_to_controller_tlast = _57;
    assign controller_to_compute_phase_1_tready = _17;
    assign controller_to_compute_phase_2_tready = _41;

endmodule
